* SPICE3 file created from RING_OSCILLATOR_0.ext - technology: sky130A

X1 VCC GND INP RING_OSCILLATOR_0

V1 VCC GND 1.8

.lib ~/open_pdks/sources/sky130-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt
.options savecurrents
.control
tran 1n 800n 790n 
*set color0=rgb:f/f/f
*set color1=rgb:0/0/0
plot  v(inp) 
.endc


.subckt RING_OSCILLATOR_0 VCC GND INP
X0 INP li_1093_1495# GND GND sky130_fd_pr__nfet_01v8 w=2.52e+06u l=150000u
X1 GND li_1093_1495# INP GND sky130_fd_pr__nfet_01v8 w=2.52e+06u l=150000u
X2 INP li_1093_1495# VCC VCC sky130_fd_pr__pfet_01v8 w=2.52e+06u l=150000u
X3 VCC li_1093_1495# INP VCC sky130_fd_pr__pfet_01v8 w=2.52e+06u l=150000u
X4 li_1093_1495# STAGE2_INV_2455088_PG0_0_0_1678382968_0/li_405_571# GND GND sky130_fd_pr__nfet_01v8 w=2.52e+06u l=150000u
X5 GND STAGE2_INV_2455088_PG0_0_0_1678382968_0/li_405_571# li_1093_1495# GND sky130_fd_pr__nfet_01v8 w=2.52e+06u l=150000u
X6 STAGE2_INV_2455088_PG0_0_0_1678382968_0/li_405_571# INP GND GND sky130_fd_pr__nfet_01v8 l=150000u
X7 GND INP STAGE2_INV_2455088_PG0_0_0_1678382968_0/li_405_571# GND sky130_fd_pr__nfet_01v8 l=150000u
X8 li_1093_1495# STAGE2_INV_2455088_PG0_0_0_1678382968_0/li_405_571# VCC VCC sky130_fd_pr__pfet_01v8 w=2.52e+06u l=150000u
X9 VCC STAGE2_INV_2455088_PG0_0_0_1678382968_0/li_405_571# li_1093_1495# VCC sky130_fd_pr__pfet_01v8 w=2.52e+06u l=150000u
X10 STAGE2_INV_2455088_PG0_0_0_1678382968_0/li_405_571# INP VCC VCC sky130_fd_pr__pfet_01v8 w=2.52e+06u l=150000u
X11 VCC INP STAGE2_INV_2455088_PG0_0_0_1678382968_0/li_405_571# VCC sky130_fd_pr__pfet_01v8 w=2.52e+06u l=150000u
C0 INP STAGE2_INV_2455088_PG0_0_0_1678382968_0/li_405_571# 0.61fF
C1 INP li_1093_1495# 0.66fF
C2 STAGE2_INV_2455088_PG0_0_0_1678382968_0/li_405_571# VCC 2.62fF
C3 VCC li_1093_1495# 2.71fF
C4 INP VCC 2.58fF
C5 STAGE2_INV_2455088_PG0_0_0_1678382968_0/li_405_571# li_1093_1495# 0.49fF
C6 INP GND 1.06fF
C7 li_1093_1495# GND 2.23fF 
C8 VCC GND 11.97fF
.ends
