* NGSPICE file created from ANALOG_0.ext - technology: sky130A

.subckt NMOS_S_25628869_X1_Y1_1677518941_1677518943 a_200_252# a_230_483# a_147_483#
X0 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_230_483# a_200_252# 0.11fF
C1 a_230_483# a_147_483# 0.74fF
C2 a_200_252# a_147_483# 0.89fF
.ends

.subckt PMOS_S_89421238_X1_Y1_1677518942_1677518943 a_200_252# a_230_399# w_0_0# VSUBS
X0 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=3.92e+06u as=8.904e+11p ps=7.78e+06u w=1.68e+06u l=150000u
X1 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
C0 a_200_252# w_0_0# 0.66fF
C1 a_200_252# a_230_399# 0.10fF
C2 a_230_399# w_0_0# 0.78fF
C3 a_230_399# VSUBS -0.03fF
C4 a_200_252# VSUBS 0.06fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt INV_21850877_PG0_0_0_1677518943 m1_54_560# li_61_1411# PMOS_S_89421238_X1_Y1_1677518942_1677518943_0/w_0_0#
+ VSUBS
XNMOS_S_25628869_X1_Y1_1677518941_1677518943_0 m1_54_560# li_61_1411# VSUBS NMOS_S_25628869_X1_Y1_1677518941_1677518943
XPMOS_S_89421238_X1_Y1_1677518942_1677518943_0 m1_54_560# li_61_1411# PMOS_S_89421238_X1_Y1_1677518942_1677518943_0/w_0_0#
+ VSUBS PMOS_S_89421238_X1_Y1_1677518942_1677518943
C0 m1_54_560# PMOS_S_89421238_X1_Y1_1677518942_1677518943_0/w_0_0# 0.29fF
C1 m1_54_560# li_61_1411# 0.17fF
C2 li_61_1411# PMOS_S_89421238_X1_Y1_1677518942_1677518943_0/w_0_0# 0.03fF
C3 li_61_1411# VSUBS 0.71fF
C4 m1_54_560# VSUBS 1.28fF
C5 PMOS_S_89421238_X1_Y1_1677518942_1677518943_0/w_0_0# VSUBS 3.02fF
.ends

.subckt PMOS_S_89421238_X1_Y1_1677518946 a_200_252# a_230_399# w_0_0# VSUBS
X0 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=3.92e+06u as=8.904e+11p ps=7.78e+06u w=1.68e+06u l=150000u
X1 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
C0 a_230_399# a_200_252# 0.10fF
C1 a_230_399# w_0_0# 0.78fF
C2 w_0_0# a_200_252# 0.66fF
C3 a_230_399# VSUBS -0.03fF
C4 a_200_252# VSUBS 0.06fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt CAP_2T_51284459_1677518944 m3_53_2692# m3_53_172# VSUBS
X0 m3_53_172# m3_53_2692# sky130_fd_pr__cap_mim_m3_1 l=10u w=10u
C0 m3_53_2692# m3_53_172# 0.83fF
C1 m3_53_172# VSUBS 0.82fF
C2 m3_53_2692# VSUBS 2.99fF
.ends

.subckt NMOS_S_25628869_X1_Y1_1677518945 a_200_252# a_230_483# a_147_483#
X0 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_200_252# a_230_483# 0.11fF
C1 a_230_483# a_147_483# 0.74fF
C2 a_200_252# a_147_483# 0.89fF
.ends

.subckt ANALOG_0 VN VP Y
XINV_21850877_PG0_0_0_1677518943_0 m3_4458_5710# Y VP VN INV_21850877_PG0_0_0_1677518943
XPMOS_S_89421238_X1_Y1_1677518946_0 Y m3_2074_2510# VP VN PMOS_S_89421238_X1_Y1_1677518946
XPMOS_S_89421238_X1_Y1_1677518946_1 m3_2074_2510# m3_4458_5710# VP VN PMOS_S_89421238_X1_Y1_1677518946
XCAP_2T_51284459_1677518944_0 Y VN VN CAP_2T_51284459_1677518944
XCAP_2T_51284459_1677518944_1 m3_4458_5710# VN VN CAP_2T_51284459_1677518944
XCAP_2T_51284459_1677518944_2 m3_2074_2510# VN VN CAP_2T_51284459_1677518944
XNMOS_S_25628869_X1_Y1_1677518945_0 m3_2074_2510# m3_4458_5710# VN NMOS_S_25628869_X1_Y1_1677518945
XNMOS_S_25628869_X1_Y1_1677518945_1 Y m3_2074_2510# VN NMOS_S_25628869_X1_Y1_1677518945
C0 m3_2074_2510# m3_4458_5710# 0.32fF
C1 m3_2074_2510# VP 7.10fF
C2 VP m3_4458_5710# 1.55fF
C3 Y m3_2074_2510# 0.90fF
C4 Y m3_4458_5710# 0.49fF
C5 Y VP 1.71fF
C6 Y VN 6.25fF
C7 m3_2074_2510# VN 6.03fF
C8 VP VN 15.82fF
C9 m3_4458_5710# VN 5.43fF
.ends



X1 VN VP Y ANALOG_0
V1 VP VN 1.8
.save i(v1)
**** begin user architecture code


.lib ~/open_pdks/sources/sky130-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt
.control
save all
tran 1u 0.001
plot v(y)
.endc

.end














