* NGSPICE file created from ANALOG_0.ext - technology: sky130A
X1 VN VP Y ANALOG_0
V1 VP VN 1.8
.save i(v1)
**** begin user architecture code


.lib ~/open_pdks/sources/sky130-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt
.control
save all
tran 10000p 4000000n
plot v(y)
.endc


.subckt PMOS_S_62253992_X5_Y1_1677862246_1677862246 a_200_252# a_230_399# w_0_0# VSUBS
X0 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.772e+12p pd=2.346e+07u as=2.352e+12p ps=1.96e+07u w=1.68e+06u l=150000u
X1 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X2 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X3 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X4 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X5 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X6 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X7 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X8 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X9 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
C0 a_200_252# a_230_399# 0.49fF
C1 a_230_399# w_0_0# 3.98fF
C2 a_200_252# w_0_0# 2.47fF
C3 a_230_399# VSUBS -0.19fF
C4 a_200_252# VSUBS 0.17fF
C5 w_0_0# VSUBS 5.49fF
.ends

.subckt NMOS_S_4459928_X5_Y1_1677862245_1677862246 a_200_252# a_230_483# a_147_483#
X0 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=1.386e+12p pd=1.338e+07u as=1.176e+12p ps=1.12e+07u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_230_483# a_200_252# 0.58fF
C1 a_230_483# a_147_483# 3.72fF
C2 a_200_252# a_147_483# 3.21fF
.ends

.subckt INV_8026114_PG0_0_0_1677862246 m1_226_1400# m1_312_560# PMOS_S_62253992_X5_Y1_1677862246_1677862246_0/w_0_0#
+ VSUBS
XPMOS_S_62253992_X5_Y1_1677862246_1677862246_0 m1_312_560# m1_226_1400# PMOS_S_62253992_X5_Y1_1677862246_1677862246_0/w_0_0#
+ VSUBS PMOS_S_62253992_X5_Y1_1677862246_1677862246
XNMOS_S_4459928_X5_Y1_1677862245_1677862246_0 m1_312_560# m1_226_1400# VSUBS NMOS_S_4459928_X5_Y1_1677862245_1677862246
C0 m1_312_560# m1_226_1400# 0.34fF
C1 m1_226_1400# PMOS_S_62253992_X5_Y1_1677862246_1677862246_0/w_0_0# 0.03fF
C2 m1_312_560# PMOS_S_62253992_X5_Y1_1677862246_1677862246_0/w_0_0# 0.36fF
C3 m1_226_1400# VSUBS 3.26fF
C4 m1_312_560# VSUBS 3.61fF
C5 PMOS_S_62253992_X5_Y1_1677862246_1677862246_0/w_0_0# VSUBS 5.63fF
.ends

.subckt PMOS_S_62253992_X5_Y1_1677862246_1677862247 a_200_252# a_230_399# w_0_0# VSUBS
X0 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.772e+12p pd=2.346e+07u as=2.352e+12p ps=1.96e+07u w=1.68e+06u l=150000u
X1 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X2 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X3 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X4 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X5 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X6 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X7 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X8 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X9 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
C0 w_0_0# a_200_252# 2.47fF
C1 w_0_0# a_230_399# 3.98fF
C2 a_230_399# a_200_252# 0.49fF
C3 a_230_399# VSUBS -0.19fF
C4 a_200_252# VSUBS 0.17fF
C5 w_0_0# VSUBS 5.49fF
.ends

.subckt NMOS_S_4459928_X5_Y1_1677862245_1677862247 a_200_252# a_230_483# a_147_483#
X0 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=1.386e+12p pd=1.338e+07u as=1.176e+12p ps=1.12e+07u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X3 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X5 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X7 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X9 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_200_252# a_230_483# 0.58fF
C1 a_230_483# a_147_483# 3.72fF
C2 a_200_252# a_147_483# 3.21fF
.ends

.subckt STAGE2_INV_31651850_PG0_0_0_1677862247 li_1093_571# m1_914_1400# m1_2032_560#
+ PMOS_S_62253992_X5_Y1_1677862246_1677862247_1/w_0_0# VSUBS
XPMOS_S_62253992_X5_Y1_1677862246_1677862247_1 m1_2032_560# li_1093_571# PMOS_S_62253992_X5_Y1_1677862246_1677862247_1/w_0_0#
+ VSUBS PMOS_S_62253992_X5_Y1_1677862246_1677862247
XPMOS_S_62253992_X5_Y1_1677862246_1677862247_0 li_1093_571# m1_914_1400# PMOS_S_62253992_X5_Y1_1677862246_1677862247_1/w_0_0#
+ VSUBS PMOS_S_62253992_X5_Y1_1677862246_1677862247
XNMOS_S_4459928_X5_Y1_1677862245_1677862247_0 li_1093_571# m1_914_1400# VSUBS NMOS_S_4459928_X5_Y1_1677862245_1677862247
XNMOS_S_4459928_X5_Y1_1677862245_1677862247_1 m1_2032_560# li_1093_571# VSUBS NMOS_S_4459928_X5_Y1_1677862245_1677862247
C0 m1_2032_560# PMOS_S_62253992_X5_Y1_1677862246_1677862247_1/w_0_0# 0.45fF
C1 li_1093_571# PMOS_S_62253992_X5_Y1_1677862246_1677862247_1/w_0_0# 1.59fF
C2 m1_914_1400# PMOS_S_62253992_X5_Y1_1677862246_1677862247_1/w_0_0# -0.00fF
C3 li_1093_571# m1_2032_560# 0.47fF
C4 m1_914_1400# m1_2032_560# 0.01fF
C5 li_1093_571# m1_914_1400# 0.07fF
C6 m1_914_1400# VSUBS 3.12fF
C7 li_1093_571# VSUBS 4.98fF
C8 PMOS_S_62253992_X5_Y1_1677862246_1677862247_1/w_0_0# VSUBS 10.48fF
C9 m1_2032_560# VSUBS 3.64fF
.ends

.subckt ANALOG_0 VN VP Y
XINV_8026114_PG0_0_0_1677862246_0 Y m2_316_1475# VP VN INV_8026114_PG0_0_0_1677862246
XSTAGE2_INV_31651850_PG0_0_0_1677862247_0 STAGE2_INV_31651850_PG0_0_0_1677862247_0/li_1093_571#
+ m2_316_1475# Y VP VN STAGE2_INV_31651850_PG0_0_0_1677862247
C0 Y STAGE2_INV_31651850_PG0_0_0_1677862247_0/li_1093_571# 0.24fF
C1 VP STAGE2_INV_31651850_PG0_0_0_1677862247_0/li_1093_571# 0.76fF
C2 m2_316_1475# Y 0.63fF
C3 m2_316_1475# VP 1.58fF
C4 Y VP 1.40fF
C5 m2_316_1475# STAGE2_INV_31651850_PG0_0_0_1677862247_0/li_1093_571# 0.47fF
C6 STAGE2_INV_31651850_PG0_0_0_1677862247_0/li_1093_571# VN 5.30fF
C7 VP VN 20.56fF
C8 Y VN 5.62fF
C9 m2_316_1475# VN 8.39fF
.ends

