magic
tech sky130A
magscale 1 2
timestamp 1676458286
<< locali >>
rect 405 1579 413 1613
rect 447 1579 455 1613
rect 405 1445 455 1579
rect 405 1411 413 1445
rect 447 1411 455 1445
<< viali >>
rect 413 1579 447 1613
rect 413 1411 447 1445
<< metal1 >>
rect 398 2462 462 2464
rect 398 2410 404 2462
rect 456 2410 462 2462
rect 398 2408 462 2410
rect 396 1613 464 1624
rect 396 1579 413 1613
rect 447 1579 464 1613
rect 396 1568 464 1579
rect 396 1445 464 1456
rect 396 1411 413 1445
rect 447 1411 464 1445
rect 396 1400 464 1411
rect 398 614 462 616
rect 398 562 404 614
rect 456 562 462 614
rect 398 560 462 562
<< via1 >>
rect 404 2410 456 2462
rect 404 562 456 614
<< metal2 >>
rect 402 2462 458 2468
rect 402 2410 404 2462
rect 456 2410 458 2462
rect 402 614 458 2410
rect 402 562 404 614
rect 456 562 458 614
rect 402 556 458 562
use NMOS_S_96839798_X1_Y1_1676446837_1676446838  NMOS_S_96839798_X1_Y1_1676446837_1676446838_0
timestamp 1676458286
transform -1 0 516 0 -1 1512
box 52 56 395 1482
use PMOS_S_36030836_X1_Y1_1676446838_1676446838  PMOS_S_36030836_X1_Y1_1676446838_1676446838_0
timestamp 1676458286
transform -1 0 516 0 1 1512
box 0 0 516 1512
<< end >>
