module analog_ring_osc(
    input in_ring,
    output rimg_adc
);

endmodule