magic
tech sky130A
magscale 1 2
timestamp 1677466831
<< locali >>
rect 405 2419 413 2453
rect 447 2419 455 2453
rect 405 2369 455 2419
rect 405 2335 413 2369
rect 447 2335 455 2369
rect 577 2335 585 2369
rect 619 2335 627 2369
rect 577 1613 627 2335
rect 405 1579 413 1613
rect 447 1579 455 1613
rect 405 1445 455 1579
rect 405 1411 413 1445
rect 447 1411 455 1445
rect 577 1579 585 1613
rect 619 1579 627 1613
rect 577 1445 627 1579
rect 577 1411 585 1445
rect 619 1411 627 1445
rect 577 1277 627 1411
rect 405 1243 413 1277
rect 447 1243 455 1277
rect 577 1243 585 1277
rect 619 1243 627 1277
rect 405 605 455 1243
rect 405 571 413 605
rect 447 571 455 605
<< viali >>
rect 413 2419 447 2453
rect 413 2335 447 2369
rect 585 2335 619 2369
rect 413 1579 447 1613
rect 413 1411 447 1445
rect 585 1579 619 1613
rect 585 1411 619 1445
rect 413 1243 447 1277
rect 585 1243 619 1277
rect 413 571 447 605
<< metal1 >>
rect 396 2453 464 2464
rect 396 2419 413 2453
rect 447 2419 464 2453
rect 396 2408 464 2419
rect 742 2462 806 2464
rect 742 2410 748 2462
rect 800 2410 806 2462
rect 742 2408 806 2410
rect 396 2369 636 2380
rect 396 2335 413 2369
rect 447 2335 585 2369
rect 619 2335 636 2369
rect 396 2324 636 2335
rect 396 1613 464 1624
rect 396 1579 413 1613
rect 447 1579 464 1613
rect 396 1568 464 1579
rect 568 1613 636 1624
rect 568 1579 585 1613
rect 619 1579 636 1613
rect 568 1568 636 1579
rect 396 1445 464 1456
rect 396 1411 413 1445
rect 447 1411 464 1445
rect 396 1400 464 1411
rect 568 1445 636 1456
rect 568 1411 585 1445
rect 619 1411 636 1445
rect 568 1400 636 1411
rect 396 1277 636 1288
rect 396 1243 413 1277
rect 447 1243 585 1277
rect 619 1243 636 1277
rect 396 1232 636 1243
rect 396 605 464 616
rect 396 571 413 605
rect 447 571 464 605
rect 396 560 464 571
rect 742 614 806 616
rect 742 562 748 614
rect 800 562 806 614
rect 742 560 806 562
<< via1 >>
rect 748 2410 800 2462
rect 748 562 800 614
<< metal2 >>
rect 746 2462 802 2468
rect 746 2410 748 2462
rect 800 2410 802 2462
rect 746 614 802 2410
rect 746 562 748 614
rect 800 562 802 614
rect 746 556 802 562
use NMOS_S_25628869_X1_Y1_1677466711_1677466713  NMOS_S_25628869_X1_Y1_1677466711_1677466713_0
timestamp 1677466831
transform -1 0 516 0 -1 1512
box 52 56 395 1482
use NMOS_S_25628869_X1_Y1_1677466711_1677466713  NMOS_S_25628869_X1_Y1_1677466711_1677466713_1
timestamp 1677466831
transform 1 0 516 0 -1 1512
box 52 56 395 1482
use PMOS_S_89421238_X1_Y1_1677466712_1677466713  PMOS_S_89421238_X1_Y1_1677466712_1677466713_0
timestamp 1677466831
transform -1 0 516 0 1 1512
box 0 0 516 1512
use PMOS_S_89421238_X1_Y1_1677466712_1677466713  PMOS_S_89421238_X1_Y1_1677466712_1677466713_1
timestamp 1677466831
transform 1 0 516 0 1 1512
box 0 0 516 1512
<< end >>
