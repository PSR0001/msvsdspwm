* NGSPICE file created from ANALOG_0.ext - technology: sky130A

.subckt PMOS_S_89421238_X1_Y1_1677407593 a_200_252# a_230_399# w_0_0# VSUBS
X0 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=3.92e+06u as=8.904e+11p ps=7.78e+06u w=1.68e+06u l=150000u
X1 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
C0 a_230_399# a_200_252# 0.10fF
C1 w_0_0# a_200_252# 0.66fF
C2 w_0_0# a_230_399# 0.78fF
C3 a_230_399# VSUBS -0.03fF
C4 a_200_252# VSUBS 0.06fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt NMOS_S_25628869_X1_Y1_1677407590_1677407590 a_200_252# a_230_483# a_147_483#
X0 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_200_252# a_230_483# 0.11fF
C1 a_230_483# a_147_483# 0.74fF
C2 a_200_252# a_147_483# 0.89fF
.ends

.subckt PMOS_S_89421238_X1_Y1_1677407591_1677407590 a_200_252# a_230_399# w_0_0# VSUBS
X0 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=3.92e+06u as=8.904e+11p ps=7.78e+06u w=1.68e+06u l=150000u
X1 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
C0 a_230_399# a_200_252# 0.10fF
C1 w_0_0# a_200_252# 0.66fF
C2 w_0_0# a_230_399# 0.78fF
C3 a_230_399# VSUBS -0.03fF
C4 a_200_252# VSUBS 0.06fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt INV_21850877_0_0_1677407590 li_405_1411# PMOS_S_89421238_X1_Y1_1677407591_1677407590_0/w_0_0#
+ m1_226_560# VSUBS
XNMOS_S_25628869_X1_Y1_1677407590_1677407590_0 m1_226_560# li_405_1411# VSUBS NMOS_S_25628869_X1_Y1_1677407590_1677407590
XPMOS_S_89421238_X1_Y1_1677407591_1677407590_0 m1_226_560# li_405_1411# PMOS_S_89421238_X1_Y1_1677407591_1677407590_0/w_0_0#
+ VSUBS PMOS_S_89421238_X1_Y1_1677407591_1677407590
C0 m1_226_560# li_405_1411# 0.14fF
C1 m1_226_560# PMOS_S_89421238_X1_Y1_1677407591_1677407590_0/w_0_0# 0.40fF
C2 PMOS_S_89421238_X1_Y1_1677407591_1677407590_0/w_0_0# li_405_1411# 0.02fF
C3 li_405_1411# VSUBS 0.68fF
C4 PMOS_S_89421238_X1_Y1_1677407591_1677407590_0/w_0_0# VSUBS 3.02fF
C5 m1_226_560# VSUBS 1.76fF
.ends

.subckt NMOS_S_25628869_X1_Y1_1677407592 a_200_252# a_230_483# a_147_483#
X0 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_200_252# a_230_483# 0.11fF
C1 a_230_483# a_147_483# 0.74fF
C2 a_200_252# a_147_483# 0.89fF
.ends

.subckt CAP_2T_9576091_1677407591 m3_53_172# m3_53_928# VSUBS
X0 m3_53_172# m3_53_928# sky130_fd_pr__cap_mim_m3_1 l=1e+06u w=1e+06u
C0 m3_53_928# m3_53_172# 0.23fF
C1 m3_53_172# VSUBS 0.30fF
C2 m3_53_928# VSUBS 0.39fF
.ends

.subckt ANALOG_0 VP Y
XPMOS_S_89421238_X1_Y1_1677407593_1 m1_430_560# m2_918_2483# VP VSUBS PMOS_S_89421238_X1_Y1_1677407593
XINV_21850877_0_0_1677407590_0 Y VP m2_918_2483# VSUBS INV_21850877_0_0_1677407590
XNMOS_S_25628869_X1_Y1_1677407592_0 m1_430_560# m2_918_2483# VSUBS NMOS_S_25628869_X1_Y1_1677407592
XNMOS_S_25628869_X1_Y1_1677407592_1 Y m1_430_560# VSUBS NMOS_S_25628869_X1_Y1_1677407592
XCAP_2T_9576091_1677407591_0 VSUBS Y VSUBS CAP_2T_9576091_1677407591
XCAP_2T_9576091_1677407591_1 VSUBS m2_918_2483# VSUBS CAP_2T_9576091_1677407591
XCAP_2T_9576091_1677407591_2 VSUBS m1_430_560# VSUBS CAP_2T_9576091_1677407591
XPMOS_S_89421238_X1_Y1_1677407593_0 Y m1_430_560# VP VSUBS PMOS_S_89421238_X1_Y1_1677407593
C0 VP Y 1.03fF
C1 m2_918_2483# VP 0.56fF
C2 VP m1_430_560# 1.59fF
C3 m2_918_2483# Y 0.25fF
C4 Y m1_430_560# 1.01fF
C5 m2_918_2483# m1_430_560# 0.51fF
C6 m1_430_560# VSUBS 2.00fF
C7 Y VSUBS 1.67fF
C8 m2_918_2483# VSUBS 2.43fF
C9 VP VSUBS 6.82fF
.ends

