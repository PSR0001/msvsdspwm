magic
tech sky130A
magscale 1 2
timestamp 1677862335
<< pwell >>
rect 215 1206 989 1482
rect 121 457 1083 677
<< nmos >>
rect 200 483 230 651
rect 286 483 316 651
rect 372 483 402 651
rect 458 483 488 651
rect 544 483 574 651
rect 630 483 660 651
rect 716 483 746 651
rect 802 483 832 651
rect 888 483 918 651
rect 974 483 1004 651
<< ndiff >>
rect 147 601 200 651
rect 147 567 155 601
rect 189 567 200 601
rect 147 533 200 567
rect 147 499 155 533
rect 189 499 200 533
rect 147 483 200 499
rect 230 601 286 651
rect 230 567 241 601
rect 275 567 286 601
rect 230 533 286 567
rect 230 499 241 533
rect 275 499 286 533
rect 230 483 286 499
rect 316 601 372 651
rect 316 567 327 601
rect 361 567 372 601
rect 316 533 372 567
rect 316 499 327 533
rect 361 499 372 533
rect 316 483 372 499
rect 402 601 458 651
rect 402 567 413 601
rect 447 567 458 601
rect 402 533 458 567
rect 402 499 413 533
rect 447 499 458 533
rect 402 483 458 499
rect 488 601 544 651
rect 488 567 499 601
rect 533 567 544 601
rect 488 533 544 567
rect 488 499 499 533
rect 533 499 544 533
rect 488 483 544 499
rect 574 601 630 651
rect 574 567 585 601
rect 619 567 630 601
rect 574 533 630 567
rect 574 499 585 533
rect 619 499 630 533
rect 574 483 630 499
rect 660 601 716 651
rect 660 567 671 601
rect 705 567 716 601
rect 660 533 716 567
rect 660 499 671 533
rect 705 499 716 533
rect 660 483 716 499
rect 746 601 802 651
rect 746 567 757 601
rect 791 567 802 601
rect 746 533 802 567
rect 746 499 757 533
rect 791 499 802 533
rect 746 483 802 499
rect 832 601 888 651
rect 832 567 843 601
rect 877 567 888 601
rect 832 533 888 567
rect 832 499 843 533
rect 877 499 888 533
rect 832 483 888 499
rect 918 601 974 651
rect 918 567 929 601
rect 963 567 974 601
rect 918 533 974 567
rect 918 499 929 533
rect 963 499 974 533
rect 918 483 974 499
rect 1004 601 1057 651
rect 1004 567 1015 601
rect 1049 567 1057 601
rect 1004 533 1057 567
rect 1004 499 1015 533
rect 1049 499 1057 533
rect 1004 483 1057 499
<< ndiffc >>
rect 155 567 189 601
rect 155 499 189 533
rect 241 567 275 601
rect 241 499 275 533
rect 327 567 361 601
rect 327 499 361 533
rect 413 567 447 601
rect 413 499 447 533
rect 499 567 533 601
rect 499 499 533 533
rect 585 567 619 601
rect 585 499 619 533
rect 671 567 705 601
rect 671 499 705 533
rect 757 567 791 601
rect 757 499 791 533
rect 843 567 877 601
rect 843 499 877 533
rect 929 567 963 601
rect 929 499 963 533
rect 1015 567 1049 601
rect 1015 499 1049 533
<< psubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
rect 413 1361 447 1456
rect 413 1232 447 1327
rect 585 1361 619 1456
rect 585 1232 619 1327
rect 757 1361 791 1456
rect 757 1232 791 1327
rect 929 1361 963 1456
rect 929 1232 963 1327
<< psubdiffcont >>
rect 241 1327 275 1361
rect 413 1327 447 1361
rect 585 1327 619 1361
rect 757 1327 791 1361
rect 929 1327 963 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 651 230 897
rect 286 651 316 897
rect 372 941 488 951
rect 372 907 413 941
rect 447 907 488 941
rect 372 897 488 907
rect 372 651 402 897
rect 458 651 488 897
rect 544 941 660 951
rect 544 907 585 941
rect 619 907 660 941
rect 544 897 660 907
rect 544 651 574 897
rect 630 651 660 897
rect 716 941 832 951
rect 716 907 757 941
rect 791 907 832 941
rect 716 897 832 907
rect 716 651 746 897
rect 802 651 832 897
rect 888 941 1004 951
rect 888 907 929 941
rect 963 907 1004 941
rect 888 897 1004 907
rect 888 651 918 897
rect 974 651 1004 897
rect 200 252 230 483
rect 286 252 316 483
rect 372 252 402 483
rect 458 252 488 483
rect 544 252 574 483
rect 630 252 660 483
rect 716 252 746 483
rect 802 252 832 483
rect 888 252 918 483
rect 974 252 1004 483
<< polycont >>
rect 241 907 275 941
rect 413 907 447 941
rect 585 907 619 941
rect 757 907 791 941
rect 929 907 963 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 405 1361 455 1445
rect 405 1327 413 1361
rect 447 1327 455 1361
rect 405 1243 455 1327
rect 577 1361 627 1445
rect 577 1327 585 1361
rect 619 1327 627 1361
rect 577 1243 627 1327
rect 749 1361 799 1445
rect 749 1327 757 1361
rect 791 1327 799 1361
rect 749 1243 799 1327
rect 921 1361 971 1445
rect 921 1327 929 1361
rect 963 1327 971 1361
rect 921 1243 971 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 405 941 455 1025
rect 405 907 413 941
rect 447 907 455 941
rect 405 823 455 907
rect 577 941 627 1025
rect 577 907 585 941
rect 619 907 627 941
rect 577 823 627 907
rect 749 941 799 1025
rect 749 907 757 941
rect 791 907 799 941
rect 749 823 799 907
rect 921 941 971 1025
rect 921 907 929 941
rect 963 907 971 941
rect 921 823 971 907
rect 147 601 197 773
rect 147 567 155 601
rect 189 567 197 601
rect 147 533 197 567
rect 147 499 155 533
rect 189 499 197 533
rect 147 185 197 499
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 601 283 773
rect 233 567 241 601
rect 275 567 283 601
rect 233 533 283 567
rect 233 499 241 533
rect 275 499 283 533
rect 233 101 283 499
rect 233 67 241 101
rect 275 67 283 101
rect 319 601 369 773
rect 319 567 327 601
rect 361 567 369 601
rect 319 533 369 567
rect 319 499 327 533
rect 361 499 369 533
rect 319 185 369 499
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
rect 405 601 455 773
rect 405 567 413 601
rect 447 567 455 601
rect 405 533 455 567
rect 405 499 413 533
rect 447 499 455 533
rect 405 101 455 499
rect 405 67 413 101
rect 447 67 455 101
rect 491 601 541 773
rect 491 567 499 601
rect 533 567 541 601
rect 491 533 541 567
rect 491 499 499 533
rect 533 499 541 533
rect 491 185 541 499
rect 491 151 499 185
rect 533 151 541 185
rect 491 67 541 151
rect 577 601 627 773
rect 577 567 585 601
rect 619 567 627 601
rect 577 533 627 567
rect 577 499 585 533
rect 619 499 627 533
rect 577 101 627 499
rect 577 67 585 101
rect 619 67 627 101
rect 663 601 713 773
rect 663 567 671 601
rect 705 567 713 601
rect 663 533 713 567
rect 663 499 671 533
rect 705 499 713 533
rect 663 185 713 499
rect 663 151 671 185
rect 705 151 713 185
rect 663 67 713 151
rect 749 601 799 773
rect 749 567 757 601
rect 791 567 799 601
rect 749 533 799 567
rect 749 499 757 533
rect 791 499 799 533
rect 749 101 799 499
rect 749 67 757 101
rect 791 67 799 101
rect 835 601 885 773
rect 835 567 843 601
rect 877 567 885 601
rect 835 533 885 567
rect 835 499 843 533
rect 877 499 885 533
rect 835 185 885 499
rect 835 151 843 185
rect 877 151 885 185
rect 835 67 885 151
rect 921 601 971 773
rect 921 567 929 601
rect 963 567 971 601
rect 921 533 971 567
rect 921 499 929 533
rect 963 499 971 533
rect 921 101 971 499
rect 921 67 929 101
rect 963 67 971 101
rect 1007 601 1057 773
rect 1007 567 1015 601
rect 1049 567 1057 601
rect 1007 533 1057 567
rect 1007 499 1015 533
rect 1049 499 1057 533
rect 1007 185 1057 499
rect 1007 151 1015 185
rect 1049 151 1057 185
rect 1007 67 1057 151
<< viali >>
rect 241 1327 275 1361
rect 413 1327 447 1361
rect 585 1327 619 1361
rect 757 1327 791 1361
rect 929 1327 963 1361
rect 241 907 275 941
rect 413 907 447 941
rect 585 907 619 941
rect 757 907 791 941
rect 929 907 963 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
rect 413 67 447 101
rect 499 151 533 185
rect 585 67 619 101
rect 671 151 705 185
rect 757 67 791 101
rect 843 151 877 185
rect 929 67 963 101
rect 1015 151 1049 185
<< metal1 >>
rect 224 1370 980 1372
rect 224 1361 662 1370
rect 224 1327 241 1361
rect 275 1327 413 1361
rect 447 1327 585 1361
rect 619 1327 662 1361
rect 224 1318 662 1327
rect 714 1361 980 1370
rect 714 1327 757 1361
rect 791 1327 929 1361
rect 963 1327 980 1361
rect 714 1318 980 1327
rect 224 1316 980 1318
rect 224 941 980 952
rect 224 907 241 941
rect 275 907 413 941
rect 447 907 585 941
rect 619 907 757 941
rect 791 907 929 941
rect 963 907 980 941
rect 224 896 980 907
rect 138 194 1066 196
rect 138 185 662 194
rect 714 185 1066 194
rect 138 151 155 185
rect 189 151 327 185
rect 361 151 499 185
rect 533 151 662 185
rect 714 151 843 185
rect 877 151 1015 185
rect 1049 151 1066 185
rect 138 142 662 151
rect 714 142 1066 151
rect 138 140 1066 142
rect 224 101 980 112
rect 224 67 241 101
rect 275 67 413 101
rect 447 67 585 101
rect 619 67 757 101
rect 791 67 929 101
rect 963 67 980 101
rect 224 56 980 67
<< via1 >>
rect 662 1318 714 1370
rect 662 185 714 194
rect 662 151 671 185
rect 671 151 705 185
rect 705 151 714 185
rect 662 142 714 151
<< metal2 >>
rect 660 1370 716 1376
rect 660 1318 662 1370
rect 714 1318 716 1370
rect 660 194 716 1318
rect 660 142 662 194
rect 714 142 716 194
rect 660 136 716 142
<< end >>
