magic
tech sky130A
magscale 1 2
timestamp 1677552377
<< error_s >>
rect 402 1083 437 1117
rect 403 1064 437 1083
rect 229 1015 287 1021
rect 229 981 241 1015
rect 229 975 287 981
rect 133 719 191 725
rect 133 685 145 719
rect 133 679 191 685
rect 422 583 437 1064
rect 456 1030 491 1064
rect 875 1030 910 1064
rect 456 583 490 1030
rect 876 1011 910 1030
rect 702 962 760 968
rect 702 928 714 962
rect 702 922 760 928
rect 606 666 664 672
rect 606 632 618 666
rect 606 626 664 632
rect 456 549 471 583
rect 895 530 910 1011
rect 929 977 964 1011
rect 929 530 963 977
rect 1175 909 1233 915
rect 1175 875 1187 909
rect 1349 892 1383 910
rect 1175 869 1233 875
rect 1349 856 1419 892
rect 1366 822 1437 856
rect 1821 822 1856 856
rect 1079 613 1137 619
rect 1079 579 1091 613
rect 1079 573 1137 579
rect 929 496 944 530
rect 1366 477 1436 822
rect 1822 803 1856 822
rect 1648 754 1706 760
rect 1648 720 1660 754
rect 1648 714 1706 720
rect 1552 560 1610 566
rect 1552 526 1564 560
rect 1552 520 1610 526
rect 1366 441 1419 477
rect 1841 424 1856 803
rect 1875 769 1910 803
rect 2294 769 2329 803
rect 1875 424 1909 769
rect 2295 750 2329 769
rect 2121 701 2179 707
rect 2121 667 2133 701
rect 2121 661 2179 667
rect 2025 507 2083 513
rect 2025 473 2037 507
rect 2025 467 2083 473
rect 1875 390 1890 424
rect 2314 371 2329 750
rect 2348 716 2383 750
rect 2348 371 2382 716
rect 2594 648 2652 654
rect 2594 614 2606 648
rect 2594 608 2652 614
rect 2498 454 2556 460
rect 2498 420 2510 454
rect 2498 414 2556 420
rect 2348 337 2363 371
<< metal1 >>
rect 0 0 200 200
rect 0 -400 200 -200
rect 0 -800 200 -600
use sky130_fd_pr__pfet_01v8_MQKFPY  XM1
timestamp 1677552377
transform 1 0 683 0 1 797
box -263 -303 263 303
use sky130_fd_pr__pfet_01v8_MQKFPY  XM2
timestamp 1677552377
transform 1 0 210 0 1 850
box -263 -303 263 303
use sky130_fd_pr__pfet_01v8_MQKFPY  XM3
timestamp 1677552377
transform 1 0 1156 0 1 744
box -263 -303 263 303
use sky130_fd_pr__nfet_01v8_MVW3GX  XM4
timestamp 1677552377
transform 1 0 1629 0 1 640
box -263 -252 263 252
use sky130_fd_pr__nfet_01v8_MVW3GX  XM5
timestamp 1677552377
transform 1 0 2102 0 1 587
box -263 -252 263 252
use sky130_fd_pr__nfet_01v8_MVW3GX  XM6
timestamp 1677552377
transform 1 0 2575 0 1 534
box -263 -252 263 252
<< labels >>
flabel metal1 0 0 200 200 0 FreeSans 256 0 0 0 VN
port 0 nsew
flabel metal1 0 -400 200 -200 0 FreeSans 256 0 0 0 VP
port 1 nsew
flabel metal1 0 -800 200 -600 0 FreeSans 256 0 0 0 Y
port 2 nsew
<< end >>
