magic
tech sky130A
magscale 1 2
timestamp 1677521559
<< checkpaint >>
rect 252 2890 2852 2914
rect 210 2872 2852 2890
rect 210 2766 3032 2872
rect 172 222 3032 2766
rect 172 122 2850 222
rect 172 116 2772 122
<< error_s >>
rect 1488 1568 1496 1624
rect 1516 1568 1524 1624
rect 1488 1400 1496 1456
rect 1516 1400 1524 1456
rect 714 928 721 1036
rect 774 868 781 986
<< locali >>
rect 577 3091 585 3125
rect 619 3091 627 3125
rect 577 2453 627 3091
rect 577 2419 585 2453
rect 619 2419 627 2453
rect 1007 2083 1015 2117
rect 1049 2083 1057 2117
rect 1007 1445 1057 2083
rect 1007 1411 1015 1445
rect 1049 1411 1057 1445
rect 1609 1579 1617 1613
rect 1651 1579 1659 1613
rect 1609 17 1659 1579
rect 1609 -17 1617 17
rect 1651 -17 1659 17
<< viali >>
rect 585 3091 619 3125
rect 585 2419 619 2453
rect 1015 2083 1049 2117
rect 1015 1411 1049 1445
rect 1617 1579 1651 1613
rect 1617 -17 1651 17
<< metal1 >>
rect 430 3974 1204 3976
rect 430 3922 576 3974
rect 628 3922 1204 3974
rect 430 3920 1204 3922
rect 54 3302 204 3304
rect 54 3250 60 3302
rect 112 3250 146 3302
rect 198 3250 204 3302
rect 54 3248 204 3250
rect 430 3125 1204 3136
rect 430 3091 585 3125
rect 619 3091 1204 3125
rect 430 3080 1204 3091
rect 570 2966 774 2968
rect 570 2914 576 2966
rect 628 2914 774 2966
rect 570 2912 774 2914
rect 568 2453 1290 2464
rect 568 2419 585 2453
rect 619 2419 1290 2453
rect 568 2408 1290 2419
rect 602 2072 774 2128
rect 946 2117 1066 2128
rect 946 2083 1015 2117
rect 1049 2083 1066 2117
rect 946 2072 1066 2083
rect 914 1622 1064 1624
rect 914 1570 920 1622
rect 972 1570 1006 1622
rect 1058 1570 1064 1622
rect 914 1568 1064 1570
rect 1550 1622 1668 1624
rect 1574 1613 1668 1622
rect 1574 1579 1617 1613
rect 1651 1579 1668 1613
rect 1574 1570 1668 1579
rect 1550 1568 1668 1570
rect 998 1454 1290 1456
rect 998 1402 1006 1454
rect 1058 1402 1290 1454
rect 998 1400 1290 1402
rect 1590 1454 1666 1456
rect 1590 1402 1608 1454
rect 1660 1402 1666 1454
rect 1590 1400 1666 1402
rect 656 1034 1322 1036
rect 656 982 662 1034
rect 714 982 1264 1034
rect 1316 982 1322 1034
rect 656 980 1322 982
rect 1600 26 1668 28
rect 1600 -26 1608 26
rect 1660 -26 1668 26
rect 1600 -28 1668 -26
<< via1 >>
rect 576 3922 628 3974
rect 60 3250 112 3302
rect 146 3250 198 3302
rect 576 2914 628 2966
rect 920 1570 972 1622
rect 1006 1570 1058 1622
rect 1550 1570 1574 1622
rect 1006 1445 1058 1454
rect 1006 1411 1015 1445
rect 1015 1411 1049 1445
rect 1049 1411 1058 1445
rect 1006 1402 1058 1411
rect 1608 1402 1660 1454
rect 662 982 714 1034
rect 1264 982 1316 1034
rect 1608 17 1660 26
rect 1608 -17 1617 17
rect 1617 -17 1651 17
rect 1651 -17 1660 17
rect 1608 -26 1660 -17
<< metal2 >>
rect 660 4060 716 4069
rect 574 3974 630 3980
rect 574 3922 576 3974
rect 628 3922 630 3974
rect 58 3302 114 3308
rect 58 3250 60 3302
rect 112 3250 114 3302
rect 58 1792 114 3250
rect 144 3302 200 3308
rect 144 3250 146 3302
rect 198 3250 200 3302
rect 144 3244 200 3250
rect 574 3304 630 3922
rect 574 2966 630 3248
rect 574 2914 576 2966
rect 628 2914 630 2966
rect 574 2908 630 2914
rect 58 1727 114 1736
rect 144 1792 200 1801
rect 144 280 200 1736
rect 316 1792 372 1801
rect 316 1727 372 1736
rect 660 1792 716 4004
rect 1434 3304 1490 3313
rect 1434 3239 1490 3248
rect 660 1727 716 1736
rect 746 1792 802 1801
rect 660 1036 716 1045
rect 660 971 716 980
rect 746 532 802 1736
rect 1606 1792 1662 1801
rect 746 467 802 476
rect 918 1622 974 1628
rect 918 1570 920 1622
rect 972 1570 974 1622
rect 144 215 200 224
rect 918 28 974 1570
rect 1004 1622 1060 1680
rect 1520 1630 1576 1680
rect 1004 1570 1006 1622
rect 1058 1570 1060 1622
rect 1004 1564 1060 1570
rect 1550 1622 1576 1630
rect 1574 1570 1576 1622
rect 1550 1564 1576 1570
rect 1004 1454 1060 1460
rect 1004 1402 1006 1454
rect 1058 1402 1060 1454
rect 1004 1288 1060 1402
rect 1606 1454 1662 1736
rect 1606 1402 1608 1454
rect 1660 1402 1662 1454
rect 1606 1396 1662 1402
rect 1520 1344 1576 1382
rect 1004 1223 1060 1232
rect 1262 1034 1318 1040
rect 1262 982 1264 1034
rect 1316 982 1318 1034
rect 1262 976 1318 982
rect 918 -37 974 -28
rect 1606 28 1662 48
rect 1606 -37 1662 -28
<< via2 >>
rect 660 4004 716 4060
rect 574 3248 630 3304
rect 58 1736 114 1792
rect 144 1736 200 1792
rect 316 1736 372 1792
rect 1434 3248 1490 3304
rect 660 1736 716 1792
rect 746 1736 802 1792
rect 660 1034 716 1036
rect 660 982 662 1034
rect 662 982 714 1034
rect 714 982 716 1034
rect 660 980 716 982
rect 1606 1736 1662 1792
rect 746 476 802 532
rect 144 224 200 280
rect 1004 1232 1060 1288
rect 918 -28 974 28
rect 1606 26 1662 28
rect 1606 -26 1608 26
rect 1608 -26 1660 26
rect 1660 -26 1662 26
rect 1606 -28 1662 -26
<< metal3 >>
rect 655 4060 721 4112
rect 655 4004 660 4060
rect 716 4004 721 4060
rect 655 3952 721 4004
rect 569 3304 635 3356
rect 569 3248 574 3304
rect 630 3248 635 3304
rect 569 3196 635 3248
rect 1429 3308 1513 3356
rect 1429 3304 1448 3308
rect 1429 3248 1434 3304
rect 1429 3244 1448 3248
rect 1512 3244 1513 3308
rect 1429 3196 1513 3244
rect -80 1796 2448 1844
rect -80 1732 -32 1796
rect 32 1792 2448 1796
rect 32 1736 58 1792
rect 114 1736 144 1792
rect 200 1736 316 1792
rect 372 1736 660 1792
rect 716 1736 746 1792
rect 802 1736 1606 1792
rect 1662 1736 2448 1792
rect 32 1732 2448 1736
rect -80 1684 2448 1732
rect 999 1288 1065 1340
rect 999 1232 1004 1288
rect 1060 1232 1065 1288
rect 999 1180 1065 1232
rect 516 1036 721 1088
rect 516 980 660 1036
rect 716 980 721 1036
rect 516 928 721 980
rect 741 532 807 584
rect 741 476 746 532
rect 802 476 807 532
rect 741 424 807 476
rect 139 280 205 332
rect 139 224 144 280
rect 200 224 205 280
rect 139 172 205 224
rect -80 32 2448 80
rect -80 28 1448 32
rect -80 -28 918 28
rect 974 -28 1448 28
rect -80 -32 1448 -28
rect 1512 28 2336 32
rect 1512 -28 1606 28
rect 1662 -28 2336 28
rect 1512 -32 2336 -28
rect 2400 -32 2448 32
rect -80 -80 2448 -32
<< via3 >>
rect 1448 3304 1512 3308
rect 1448 3248 1490 3304
rect 1490 3248 1512 3304
rect 1448 3244 1512 3248
rect -32 1732 32 1796
rect 1448 -32 1512 32
rect 2336 -32 2400 32
<< metal4 >>
rect -118 1796 118 3646
rect -118 1732 -32 1796
rect 32 1732 118 1796
rect -118 -118 118 1732
rect 1362 3308 1598 3309
rect 1362 3244 1448 3308
rect 1512 3244 1598 3308
rect 1362 1512 1598 3244
rect 1362 1506 1510 1512
rect 1362 1376 1432 1506
rect 1590 1382 1598 1512
rect 1512 1376 1598 1382
rect 1362 32 1598 1376
rect 1362 -32 1448 32
rect 1512 -32 1598 32
rect 1362 -33 1598 -32
rect 2250 32 2486 3646
rect 2250 -32 2336 32
rect 2400 -32 2486 32
rect 2250 -118 2486 -32
use CAP_2T_9576091_1677518467  CAP_2T_9576091_1677518467_0
timestamp 1677521313
transform 1 0 602 0 1 252
box 53 166 463 1088
use CAP_2T_9576091_1677518467  CAP_2T_9576091_1677518467_1
timestamp 1677521313
transform -1 0 602 0 1 0
box 53 166 463 1088
use CAP_2T_9576091_1677518467  CAP_2T_9576091_1677518467_2
timestamp 1677521313
transform 1 0 516 0 -1 4284
box 53 166 463 1088
use INV_21850877_PG0_0_0_1677518466  INV_21850877_PG0_0_0_1677518466_0
timestamp 1677521313
transform 1 0 1204 0 1 0
box 0 30 516 3024
use NMOS_S_25628869_X1_Y1_1677518468  NMOS_S_25628869_X1_Y1_1677518468_0
timestamp 1677521313
transform -1 0 516 0 1 3024
box 52 56 395 1482
use NMOS_S_25628869_X1_Y1_1677518468  NMOS_S_25628869_X1_Y1_1677518468_1
timestamp 1677521313
transform -1 0 688 0 -1 3024
box 52 56 395 1482
use PMOS_S_89421238_X1_Y1_1677518469  PMOS_S_89421238_X1_Y1_1677518469_0
timestamp 1677521313
transform 1 0 688 0 -1 3024
box 0 0 516 1512
use PMOS_S_89421238_X1_Y1_1677518469  PMOS_S_89421238_X1_Y1_1677518469_1
timestamp 1677521313
transform 1 0 1118 0 1 3024
box 0 0 516 1512
<< labels >>
flabel metal3 s 860 1260 860 1260 0 FreeSerif 0 0 0 0 Y
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal2 s 688 2898 688 2898 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 2646 0 2646 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal3 s 1471 3276 1471 3276 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 2368 2646 2368 2646 0 FreeSerif 0 0 0 0 VP
<< end >>
