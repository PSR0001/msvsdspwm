module analog_1bit_adc(
    input in_bias,
    input in_inn,
    output out_adc
);

(*I do not know how to write @@ codes EX: @@ @no a_buffer_0 (.A(lc_0), .nbout(lc_out)); *)

endmodule