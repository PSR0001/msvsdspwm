magic
tech sky130A
magscale 1 2
timestamp 1677522882
<< locali >>
rect 1695 5947 1703 5981
rect 1737 5947 1745 5981
rect 1695 5477 1745 5947
rect 1179 5443 1187 5477
rect 1221 5443 1229 5477
rect 1695 5443 1703 5477
rect 1737 5443 1745 5477
rect 1179 3965 1229 5443
rect 1695 4519 1703 4553
rect 1737 4519 1745 4553
rect 1695 4469 1745 4519
rect 1695 4435 1703 4469
rect 1737 4435 1745 4469
rect 1179 3931 1187 3965
rect 1221 3931 1229 3965
rect 1867 3965 1917 4452
rect 1867 3931 1875 3965
rect 1909 3931 1917 3965
<< viali >>
rect 1703 5947 1737 5981
rect 1187 5443 1221 5477
rect 1703 5443 1737 5477
rect 1703 4519 1737 4553
rect 1703 4435 1737 4469
rect 1187 3931 1221 3965
rect 1875 3931 1909 3965
<< metal1 >>
rect 1686 5981 1754 5992
rect 1686 5947 1703 5981
rect 1737 5947 1754 5981
rect 1686 5936 1754 5947
rect 1170 5477 1238 5488
rect 1170 5443 1187 5477
rect 1221 5443 1238 5477
rect 1170 5432 1238 5443
rect 1686 5477 1892 5488
rect 1686 5443 1703 5477
rect 1737 5443 1892 5477
rect 1686 5432 1892 5443
rect 2064 5486 2440 5488
rect 2064 5434 2382 5486
rect 2434 5434 2440 5486
rect 2064 5432 2440 5434
rect 2032 5318 2526 5320
rect 2032 5266 2038 5318
rect 2090 5266 2468 5318
rect 2520 5266 2526 5318
rect 2032 5264 2526 5266
rect 1516 5150 1580 5152
rect 1516 5098 1522 5150
rect 1574 5098 1580 5150
rect 1516 5096 1580 5098
rect 1204 4646 1580 4648
rect 1204 4594 1522 4646
rect 1574 4594 1580 4646
rect 1204 4592 1580 4594
rect 2186 4646 2268 4648
rect 2186 4594 2210 4646
rect 2262 4594 2268 4646
rect 2186 4592 2268 4594
rect 1686 4562 1924 4564
rect 1686 4553 1866 4562
rect 1686 4519 1703 4553
rect 1737 4519 1866 4553
rect 1686 4510 1866 4519
rect 1918 4510 1924 4562
rect 1686 4508 1924 4510
rect 828 4478 978 4480
rect 828 4426 834 4478
rect 886 4426 920 4478
rect 972 4426 978 4478
rect 828 4424 978 4426
rect 1686 4469 1754 4480
rect 1686 4435 1703 4469
rect 1737 4435 1754 4469
rect 1686 4424 1754 4435
rect 1344 4310 1494 4312
rect 1344 4258 1350 4310
rect 1402 4258 1436 4310
rect 1488 4258 1494 4310
rect 1344 4256 1494 4258
rect 1774 4310 2182 4312
rect 1774 4258 1780 4310
rect 1832 4258 2124 4310
rect 2176 4258 2182 4310
rect 1774 4256 2182 4258
rect 1170 3974 2440 3976
rect 1170 3965 2382 3974
rect 1170 3931 1187 3965
rect 1221 3931 1875 3965
rect 1909 3931 2382 3965
rect 1170 3922 2382 3931
rect 2434 3922 2440 3974
rect 1170 3920 2440 3922
rect 1000 3134 1064 3136
rect 1000 3082 1006 3134
rect 1058 3082 1064 3134
rect 1000 3080 1064 3082
rect 1270 3014 1330 3920
rect 1516 3638 1580 3640
rect 1516 3586 1522 3638
rect 1574 3586 1580 3638
rect 1516 3584 1580 3586
rect 1270 2942 4542 3014
rect 1946 2630 2440 2632
rect 1946 2578 1952 2630
rect 2004 2578 2382 2630
rect 2434 2578 2440 2630
rect 1946 2576 2440 2578
<< via1 >>
rect 2382 5434 2434 5486
rect 2038 5266 2090 5318
rect 2468 5266 2520 5318
rect 1522 5098 1574 5150
rect 1522 4594 1574 4646
rect 2210 4594 2262 4646
rect 1866 4510 1918 4562
rect 834 4426 886 4478
rect 920 4426 972 4478
rect 1350 4258 1402 4310
rect 1436 4258 1488 4310
rect 1780 4258 1832 4310
rect 2124 4258 2176 4310
rect 2382 3922 2434 3974
rect 1006 3082 1058 3134
rect 1522 3586 1574 3638
rect 1952 2578 2004 2630
rect 2382 2578 2434 2630
<< metal2 >>
rect 2380 5824 2436 5833
rect 2380 5486 2436 5768
rect 2380 5434 2382 5486
rect 2434 5434 2436 5486
rect 2380 5428 2436 5434
rect 58 5320 114 5329
rect 58 280 114 5264
rect 832 5320 888 5329
rect 832 4478 888 5264
rect 1348 5320 1404 5329
rect 918 4816 974 4825
rect 918 4751 974 4760
rect 832 4426 834 4478
rect 886 4426 888 4478
rect 832 4420 888 4426
rect 918 4478 974 4484
rect 918 4426 920 4478
rect 972 4426 974 4478
rect 918 4368 974 4426
rect 1348 4310 1404 5264
rect 1778 5320 1834 5329
rect 1520 5150 1576 5156
rect 1520 5098 1522 5150
rect 1574 5098 1576 5150
rect 1434 4816 1490 4825
rect 1434 4751 1490 4760
rect 1520 4646 1576 5098
rect 1520 4594 1522 4646
rect 1574 4594 1576 4646
rect 1348 4258 1350 4310
rect 1402 4258 1404 4310
rect 1348 4252 1404 4258
rect 1434 4310 1490 4316
rect 1434 4258 1436 4310
rect 1488 4258 1490 4310
rect 1434 4252 1490 4258
rect 1520 3638 1576 4594
rect 1778 4310 1834 5264
rect 1950 5320 2006 5329
rect 1864 4562 1920 4568
rect 1864 4510 1866 4562
rect 1918 4510 1920 4562
rect 1864 4504 1920 4510
rect 1778 4258 1780 4310
rect 1832 4258 1834 4310
rect 1778 4252 1834 4258
rect 1520 3586 1522 3638
rect 1574 3586 1576 3638
rect 1004 3134 1060 3140
rect 1004 3082 1006 3134
rect 1058 3082 1060 3134
rect 1004 2800 1060 3082
rect 1004 2735 1060 2744
rect 1520 2800 1576 3586
rect 1520 2735 1576 2744
rect 1950 2630 2006 5264
rect 2036 5320 2092 5329
rect 2036 5255 2092 5264
rect 2466 5318 2522 5324
rect 2466 5266 2468 5318
rect 2520 5266 2522 5318
rect 2124 4678 2264 4730
rect 2208 4646 2264 4678
rect 2208 4594 2210 4646
rect 2262 4594 2264 4646
rect 2122 4310 2178 4316
rect 2122 4258 2124 4310
rect 2176 4258 2178 4310
rect 2122 4252 2178 4258
rect 1950 2578 1952 2630
rect 2004 2578 2006 2630
rect 1950 2572 2006 2578
rect 58 215 114 224
rect 2208 28 2264 4594
rect 2380 3974 2436 3980
rect 2380 3922 2382 3974
rect 2434 3922 2436 3974
rect 2380 2800 2436 3922
rect 2466 3304 2522 5266
rect 2466 3239 2522 3248
rect 2380 2735 2436 2744
rect 2380 2630 2436 2636
rect 2380 2578 2382 2630
rect 2434 2578 2436 2630
rect 2380 280 2436 2578
rect 2380 215 2436 224
rect 2208 -37 2264 -28
<< via2 >>
rect 2380 5768 2436 5824
rect 58 5264 114 5320
rect 832 5264 888 5320
rect 1348 5264 1404 5320
rect 918 4760 974 4816
rect 1778 5264 1834 5320
rect 1434 4760 1490 4816
rect 1950 5264 2006 5320
rect 1004 2744 1060 2800
rect 1520 2744 1576 2800
rect 2036 5318 2092 5320
rect 2036 5266 2038 5318
rect 2038 5266 2090 5318
rect 2090 5266 2092 5318
rect 2036 5264 2092 5266
rect 58 224 114 280
rect 2466 3248 2522 3304
rect 2380 2744 2436 2800
rect 2380 224 2436 280
rect 2208 -28 2264 28
<< metal3 >>
rect -86 6258 4572 6264
rect -90 6076 4572 6258
rect -90 5372 98 6076
rect 2375 5824 2441 5876
rect 2375 5768 2380 5824
rect 2436 5768 2441 5824
rect 2375 5716 2441 5768
rect 4458 5710 4548 5874
rect -90 5320 2144 5372
rect -90 5264 58 5320
rect 114 5264 832 5320
rect 888 5264 1348 5320
rect 1404 5264 1778 5320
rect 1834 5264 1950 5320
rect 2006 5264 2036 5320
rect 2092 5264 2144 5320
rect -90 5212 2144 5264
rect 855 4820 979 4868
rect 855 4756 856 4820
rect 920 4816 979 4820
rect 974 4760 979 4816
rect 920 4756 979 4760
rect 855 4708 979 4756
rect 1429 4820 1513 4868
rect 1429 4816 1448 4820
rect 1429 4760 1434 4816
rect 1429 4756 1448 4760
rect 1512 4756 1513 4820
rect 1429 4708 1513 4756
rect 2461 3304 2527 3356
rect 2461 3248 2466 3304
rect 2522 3248 2527 3304
rect 2461 3196 2527 3248
rect 999 2800 1065 2852
rect 999 2744 1004 2800
rect 1060 2744 1065 2800
rect 999 2692 1065 2744
rect 1515 2800 1581 2852
rect 1515 2744 1520 2800
rect 1576 2744 1581 2800
rect 2375 2800 2441 2852
rect 1515 2692 1581 2744
rect 2074 2510 2158 2760
rect 2375 2744 2380 2800
rect 2436 2744 2441 2800
rect 2375 2692 2441 2744
rect 4466 2664 4554 2850
rect 53 280 119 332
rect 53 224 58 280
rect 114 224 119 280
rect 53 172 119 224
rect 2375 280 2441 332
rect 2375 224 2380 280
rect 2436 224 2441 280
rect 2375 172 2441 224
rect -88 32 4564 94
rect -88 -32 856 32
rect 920 -32 1448 32
rect 1512 28 4564 32
rect 1512 -28 2208 28
rect 2264 -28 4564 28
rect 1512 -32 4564 -28
rect -88 -82 4564 -32
<< via3 >>
rect 856 4816 920 4820
rect 856 4760 918 4816
rect 918 4760 920 4816
rect 856 4756 920 4760
rect 1448 4816 1512 4820
rect 1448 4760 1490 4816
rect 1490 4760 1512 4816
rect 1448 4756 1512 4760
rect 856 -32 920 32
rect 1448 -32 1512 32
<< metal4 >>
rect 770 4820 1006 4821
rect 770 4756 856 4820
rect 920 4756 1006 4820
rect 770 32 1006 4756
rect 770 -32 856 32
rect 920 -32 1006 32
rect 770 -33 1006 -32
rect 1362 4820 1598 4821
rect 1362 4756 1448 4820
rect 1512 4756 1598 4820
rect 1362 32 1598 4756
rect 1362 -32 1448 32
rect 1512 -32 1598 32
rect 1362 -33 1598 -32
use CAP_2T_51284459_1677518944  CAP_2T_51284459_1677518944_0
timestamp 1677519681
transform 1 0 2322 0 1 0
box 53 166 2232 2852
use CAP_2T_51284459_1677518944  CAP_2T_51284459_1677518944_1
timestamp 1677519681
transform 1 0 2322 0 1 3024
box 53 166 2232 2852
use CAP_2T_51284459_1677518944  CAP_2T_51284459_1677518944_2
timestamp 1677519681
transform 1 0 0 0 1 0
box 53 166 2232 2852
use INV_21850877_PG0_0_0_1677518943  INV_21850877_PG0_0_0_1677518943_0
timestamp 1677519681
transform 1 0 1806 0 1 3024
box 0 30 516 3024
use NMOS_S_25628869_X1_Y1_1677518945  NMOS_S_25628869_X1_Y1_1677518945_0
timestamp 1677519681
transform -1 0 1806 0 -1 4536
box 52 56 395 1482
use NMOS_S_25628869_X1_Y1_1677518945  NMOS_S_25628869_X1_Y1_1677518945_1
timestamp 1677519681
transform -1 0 1290 0 1 3024
box 52 56 395 1482
use PMOS_S_89421238_X1_Y1_1677518946  PMOS_S_89421238_X1_Y1_1677518946_0
timestamp 1677519681
transform -1 0 1290 0 1 4536
box 0 0 516 1512
use PMOS_S_89421238_X1_Y1_1677518946  PMOS_S_89421238_X1_Y1_1677518946_1
timestamp 1677519681
transform -1 0 1806 0 -1 6048
box 0 0 516 1512
<< labels >>
flabel metal3 s 1471 4788 1471 4788 0 FreeSerif 0 0 0 0 VP
rlabel metal3 486 26 486 26 1 VP
port 2 n
rlabel locali 1204 4128 1204 4128 1 Y
port 3 n
rlabel metal3 -12 6156 -12 6156 1 VN
port 1 n
<< end >>
