* SPICE3 file created from COMPARATOR_0.ext - technology: sky130A

X1 OUT VCC GND INP INN BIAS COMPARATOR_0

V2 VCC GND 1.8
V3 INN GND 1
V4 INP GND sine(0 1.8 100000000)
V1 BIAS GND 0.9

.lib ~/open_pdks/sources/sky130-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt
*.options savecurrents
.control
tran 0.1n 100n
plot v(out) v(inp)
.endc

.subckt COMPARATOR_0 OUT VCC GND INP INN BIAS
X0 m1_828_1316# INP m1_430_1652# GND sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=1.1256e+12p ps=1.108e+07u w=840000u l=150000u
X1 m1_430_1652# INP m1_828_1316# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 li_491_1495# INN m1_430_1652# GND sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=0p ps=0u w=840000u l=150000u
X3 m1_430_1652# INN li_491_1495# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X4 li_491_1495# li_491_1495# VCC VCC sky130_fd_pr__pfet_01v8 ad=2.352e+11p pd=2.24e+06u as=2.016e+12p ps=1.992e+07u w=840000u l=150000u
X5 VCC li_491_1495# li_491_1495# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X6 m1_828_1316# li_491_1495# VCC VCC sky130_fd_pr__pfet_01v8 ad=2.352e+11p pd=2.24e+06u as=0p ps=0u w=840000u l=150000u
X7 VCC li_491_1495# m1_828_1316# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X8 li_2125_1411# STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# GND GND sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=1.7808e+12p ps=1.768e+07u w=840000u l=150000u
X9 GND STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# li_2125_1411# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X10 STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# m1_828_1316# GND GND sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=0p ps=0u w=840000u l=150000u
X11 GND m1_828_1316# STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X12 li_2125_1411# STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# VCC VCC sky130_fd_pr__pfet_01v8 ad=2.352e+11p pd=2.24e+06u as=0p ps=0u w=840000u l=150000u
X13 VCC STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# li_2125_1411# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X14 STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# m1_828_1316# VCC VCC sky130_fd_pr__pfet_01v8 ad=2.352e+11p pd=2.24e+06u as=0p ps=0u w=840000u l=150000u
X15 VCC m1_828_1316# STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X16 m1_430_1652# BIAS GND GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X17 GND BIAS m1_430_1652# GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X18 OUT li_2125_1411# GND GND sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=0p ps=0u w=840000u l=150000u
X19 GND li_2125_1411# OUT GND sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X20 OUT li_2125_1411# VCC VCC sky130_fd_pr__pfet_01v8 ad=2.352e+11p pd=2.24e+06u as=0p ps=0u w=840000u l=150000u
X21 VCC li_2125_1411# OUT VCC sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 INN li_2125_1411# 0.00fF
C1 OUT li_2125_1411# 0.66fF
C2 STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# INP 0.00fF
C3 STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# m1_430_1652# 0.00fF
C4 STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# li_491_1495# 0.01fF
C5 li_2125_1411# VCC 2.93fF
C6 BIAS m1_430_1652# 0.11fF
C7 m1_828_1316# li_2125_1411# 0.03fF
C8 BIAS li_491_1495# 0.05fF
C9 INN STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# 0.00fF
C10 STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# OUT 0.00fF
C11 INN BIAS 0.00fF
C12 m1_430_1652# INP 0.12fF
C13 li_491_1495# INP 0.00fF
C14 STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# VCC 2.60fF
C15 m1_430_1652# li_491_1495# 1.01fF
C16 STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# m1_828_1316# 0.71fF
C17 INN INP 0.04fF
C18 OUT INP 0.00fF
C19 BIAS VCC 0.08fF
C20 BIAS m1_828_1316# 0.00fF
C21 INN m1_430_1652# 0.13fF
C22 OUT m1_430_1652# 0.00fF
C23 INN li_491_1495# 0.11fF
C24 OUT li_491_1495# 0.00fF
C25 VCC INP 0.04fF
C26 m1_828_1316# INP 0.15fF
C27 m1_430_1652# VCC 0.17fF
C28 STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# li_2125_1411# 0.43fF
C29 m1_828_1316# m1_430_1652# 0.68fF
C30 VCC li_491_1495# 2.61fF
C31 m1_828_1316# li_491_1495# 0.40fF
C32 INN VCC 0.00fF
C33 OUT VCC 0.95fF
C34 INN m1_828_1316# 0.00fF
C35 m1_828_1316# OUT 0.00fF
C36 li_2125_1411# INP 0.00fF
C37 m1_430_1652# li_2125_1411# 0.00fF
C38 STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# BIAS 0.00fF
C39 m1_828_1316# VCC 3.18fF
C40 li_2125_1411# li_491_1495# 0.00fF
C41 OUT GND 0.66fF
C42 m1_430_1652# GND 1.35fF 
C43 BIAS GND 0.85fF
C44 STAGE2_INV_89790208_PG0_0_0_1678373050_0/li_405_571# GND 1.23fF 
C45 m1_828_1316# GND 0.80fF 
C46 li_2125_1411# GND 1.63fF 
C47 VCC GND 15.92fF
C48 li_491_1495# GND 0.05fF 
C49 INN GND 0.82fF
C50 INP GND 0.75fF
.ends
