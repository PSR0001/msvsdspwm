* NGSPICE file created from FUNCTION_SKY130_0.ext - technology: sky130A

.subckt NMOS_S_96839798_X1_Y1_1676446840 a_147_525# a_200_252# a_230_525#
X0 a_230_525# a_200_252# a_147_525# a_147_525# sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X1 a_147_525# a_200_252# a_230_525# a_147_525# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_200_252# a_230_525# 0.12fF
C1 a_230_525# a_147_525# 0.73fF
C2 a_200_252# a_147_525# 0.97fF
.ends

.subckt PMOS_S_36030836_X1_Y1_1676446841 a_200_252# a_230_483# w_0_0# VSUBS
X0 a_230_483# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 w_0_0# a_200_252# a_230_483# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 w_0_0# a_200_252# 0.80fF
C1 a_200_252# a_230_483# 0.11fF
C2 w_0_0# a_230_483# 0.78fF
C3 a_230_483# VSUBS -0.04fF
C4 a_200_252# VSUBS 0.09fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt NMOS_S_96839798_X1_Y1_1676446837_1676446838 a_147_525# a_200_252# a_230_525#
X0 a_230_525# a_200_252# a_147_525# a_147_525# sky130_fd_pr__nfet_01v8 ad=1.176e+11p pd=1.4e+06u as=2.226e+11p ps=2.74e+06u w=420000u l=150000u
X1 a_147_525# a_200_252# a_230_525# a_147_525# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=420000u l=150000u
C0 a_200_252# a_230_525# 0.12fF
C1 a_230_525# a_147_525# 0.73fF
C2 a_200_252# a_147_525# 0.97fF
.ends

.subckt PMOS_S_36030836_X1_Y1_1676446838_1676446838 a_200_252# a_230_483# w_0_0# VSUBS
X0 a_230_483# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 w_0_0# a_200_252# a_230_483# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 w_0_0# a_200_252# 0.80fF
C1 a_200_252# a_230_483# 0.11fF
C2 w_0_0# a_230_483# 0.78fF
C3 a_230_483# VSUBS -0.04fF
C4 a_200_252# VSUBS 0.09fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt INV_6743645_0_0_1676446838 li_405_1411# PMOS_S_36030836_X1_Y1_1676446838_1676446838_0/w_0_0#
+ m1_398_560# VSUBS
XNMOS_S_96839798_X1_Y1_1676446837_1676446838_0 VSUBS m1_398_560# li_405_1411# NMOS_S_96839798_X1_Y1_1676446837_1676446838
XPMOS_S_36030836_X1_Y1_1676446838_1676446838_0 m1_398_560# li_405_1411# PMOS_S_36030836_X1_Y1_1676446838_1676446838_0/w_0_0#
+ VSUBS PMOS_S_36030836_X1_Y1_1676446838_1676446838
C0 PMOS_S_36030836_X1_Y1_1676446838_1676446838_0/w_0_0# li_405_1411# 0.06fF
C1 m1_398_560# PMOS_S_36030836_X1_Y1_1676446838_1676446838_0/w_0_0# 0.29fF
C2 m1_398_560# li_405_1411# 0.15fF
C3 li_405_1411# VSUBS 0.67fF
C4 m1_398_560# VSUBS 1.63fF
C5 PMOS_S_36030836_X1_Y1_1676446838_1676446838_0/w_0_0# VSUBS 3.02fF
.ends

.subckt DP_PMOS_90543401_X1_Y1_1676446839 a_372_252# a_200_252# a_230_483# a_402_483#
+ w_0_0# VSUBS
X0 a_230_483# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.352e+11p pd=2.24e+06u as=6.804e+11p ps=6.66e+06u w=840000u l=150000u
X1 w_0_0# a_200_252# a_230_483# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
X2 a_402_483# a_372_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=2.352e+11p pd=2.24e+06u as=0p ps=0u w=840000u l=150000u
X3 w_0_0# a_372_252# a_402_483# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_402_483# a_200_252# 0.01fF
C1 a_372_252# a_402_483# 0.12fF
C2 a_372_252# a_200_252# 0.26fF
C3 a_402_483# w_0_0# 0.91fF
C4 w_0_0# a_200_252# 0.68fF
C5 a_372_252# w_0_0# 0.69fF
C6 a_230_483# a_402_483# 0.06fF
C7 a_230_483# a_200_252# 0.12fF
C8 a_230_483# w_0_0# 0.72fF
C9 a_402_483# VSUBS -0.07fF
C10 a_230_483# VSUBS -0.11fF
C11 a_372_252# VSUBS 0.06fF
C12 a_200_252# VSUBS 0.01fF
C13 w_0_0# VSUBS 3.45fF
.ends

.subckt FUNCTION_SKY130_0
XNMOS_S_96839798_X1_Y1_1676446840_0 VSS m1_1806_2408# Y NMOS_S_96839798_X1_Y1_1676446840
XNMOS_S_96839798_X1_Y1_1676446840_1 VSS m1_1978_560# Y NMOS_S_96839798_X1_Y1_1676446840
XNMOS_S_96839798_X1_Y1_1676446840_2 VSS F VSS NMOS_S_96839798_X1_Y1_1676446840
XNMOS_S_96839798_X1_Y1_1676446840_3 VSS D VSS NMOS_S_96839798_X1_Y1_1676446840
XNMOS_S_96839798_X1_Y1_1676446840_4 VSS B VSS NMOS_S_96839798_X1_Y1_1676446840
XPMOS_S_36030836_X1_Y1_1676446841_0 m1_2838_2408# m1_312_224# VDD VSS PMOS_S_36030836_X1_Y1_1676446841
XPMOS_S_36030836_X1_Y1_1676446841_1 C m1_312_224# VDD VSS PMOS_S_36030836_X1_Y1_1676446841
XPMOS_S_36030836_X1_Y1_1676446841_2 m1_946_560# Y m1_312_224# VSS PMOS_S_36030836_X1_Y1_1676446841
XINV_6743645_0_0_1676446838_0 Y m1_312_224# E VSS INV_6743645_0_0_1676446838
XDP_PMOS_90543401_X1_Y1_1676446839_0 li_2813_487# m1_1978_560# VDD VDD VDD VSS DP_PMOS_90543401_X1_Y1_1676446839
C0 F E 0.04fF
C1 m1_312_224# m1_1978_560# 0.00fF
C2 B D 0.00fF
C3 Y m1_312_224# 0.66fF
C4 li_2813_487# VDD 0.01fF
C5 D VDD 0.16fF
C6 Y C 0.00fF
C7 C m1_312_224# 0.01fF
C8 B m1_312_224# 0.00fF
C9 Y F 0.00fF
C10 A Y 0.01fF
C11 m1_2838_2408# m1_1806_2408# 0.00fF
C12 F m1_312_224# 0.27fF
C13 A m1_312_224# 0.00fF
C14 m1_946_560# m1_1978_560# 0.00fF
C15 Y VDD 0.07fF
C16 Y m1_946_560# 0.00fF
C17 m1_312_224# VDD 1.60fF
C18 m1_946_560# m1_312_224# 0.00fF
C19 li_2813_487# m1_1978_560# 0.00fF
C20 A C 0.00fF
C21 Y E 0.04fF
C22 E m1_312_224# 0.05fF
C23 li_2813_487# m1_312_224# 0.00fF
C24 C VDD 0.25fF
C25 D m1_312_224# 0.00fF
C26 B F 0.00fF
C27 B A 0.00fF
C28 A F 0.04fF
C29 C E 0.01fF
C30 B VDD 0.26fF
C31 Y m1_1806_2408# 0.00fF
C32 D C 0.04fF
C33 F VDD 0.00fF
C34 A VDD 0.18fF
C35 m1_312_224# m1_1806_2408# 0.00fF
C36 A VSS 0.08fF $ **FLOATING
C37 VDD VSS 9.82fF
C38 li_2813_487# VSS 0.30fF
C39 m1_1978_560# VSS 1.08fF
C40 Y VSS 2.85fF
C41 E VSS 1.26fF
C42 m1_312_224# VSS 4.55fF
C43 m1_946_560# VSS 0.17fF
C44 C VSS -0.44fF
C45 m1_2838_2408# VSS 0.17fF
C46 B VSS 0.52fF
C47 D VSS 0.61fF
C48 F VSS 0.43fF
C49 m1_1806_2408# VSS 1.05fF
.ends

