* NGSPICE file created from ANALOG_0.ext - technology: sky130A

.subckt NMOS_S_25628869_X1_Y1_1677466711_1677466713 a_200_252# a_230_483# a_147_483#
X0 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_230_483# a_200_252# 0.11fF
C1 a_230_483# a_147_483# 0.74fF
C2 a_200_252# a_147_483# 0.89fF
.ends

.subckt PMOS_S_89421238_X1_Y1_1677466712_1677466713 a_200_252# a_230_399# w_0_0# VSUBS
X0 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=3.92e+06u as=8.904e+11p ps=7.78e+06u w=1.68e+06u l=150000u
X1 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
C0 a_230_399# w_0_0# 0.78fF
C1 a_200_252# w_0_0# 0.66fF
C2 a_230_399# a_200_252# 0.10fF
C3 a_230_399# VSUBS -0.03fF
C4 a_200_252# VSUBS 0.06fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt STAGE2_INV_27873531_PG0_0_0_1677466713 li_405_1411# li_405_571# PMOS_S_89421238_X1_Y1_1677466712_1677466713_1/w_0_0#
+ m1_742_560# VSUBS
XNMOS_S_25628869_X1_Y1_1677466711_1677466713_0 li_405_571# li_405_1411# VSUBS NMOS_S_25628869_X1_Y1_1677466711_1677466713
XNMOS_S_25628869_X1_Y1_1677466711_1677466713_1 m1_742_560# li_405_571# VSUBS NMOS_S_25628869_X1_Y1_1677466711_1677466713
XPMOS_S_89421238_X1_Y1_1677466712_1677466713_0 li_405_571# li_405_1411# PMOS_S_89421238_X1_Y1_1677466712_1677466713_1/w_0_0#
+ VSUBS PMOS_S_89421238_X1_Y1_1677466712_1677466713
XPMOS_S_89421238_X1_Y1_1677466712_1677466713_1 m1_742_560# li_405_571# PMOS_S_89421238_X1_Y1_1677466712_1677466713_1/w_0_0#
+ VSUBS PMOS_S_89421238_X1_Y1_1677466712_1677466713
C0 m1_742_560# li_405_571# 0.38fF
C1 li_405_1411# PMOS_S_89421238_X1_Y1_1677466712_1677466713_1/w_0_0# 0.10fF
C2 m1_742_560# PMOS_S_89421238_X1_Y1_1677466712_1677466713_1/w_0_0# 0.71fF
C3 m1_742_560# li_405_1411# 0.02fF
C4 li_405_571# PMOS_S_89421238_X1_Y1_1677466712_1677466713_1/w_0_0# 0.92fF
C5 li_405_571# li_405_1411# 0.11fF
C6 li_405_571# VSUBS 0.90fF
C7 m1_742_560# VSUBS 0.93fF
C8 li_405_1411# VSUBS 0.59fF
C9 PMOS_S_89421238_X1_Y1_1677466712_1677466713_1/w_0_0# VSUBS 5.04fF
.ends

.subckt PMOS_S_89421238_X1_Y1_1677466712_1677466712 a_200_252# a_230_399# w_0_0# VSUBS
X0 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=3.92e+06u as=8.904e+11p ps=7.78e+06u w=1.68e+06u l=150000u
X1 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
C0 w_0_0# a_230_399# 0.78fF
C1 a_230_399# a_200_252# 0.10fF
C2 w_0_0# a_200_252# 0.66fF
C3 a_230_399# VSUBS -0.03fF
C4 a_200_252# VSUBS 0.06fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt NMOS_S_25628869_X1_Y1_1677466711_1677466712 a_200_252# a_230_483# a_147_483#
X0 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_200_252# a_230_483# 0.11fF
C1 a_230_483# a_147_483# 0.74fF
C2 a_200_252# a_147_483# 0.89fF
.ends

.subckt INV_21850877_PG0_0_0_1677466712 PMOS_S_89421238_X1_Y1_1677466712_1677466712_0/w_0_0#
+ li_61_1411# m1_226_560# VSUBS
XPMOS_S_89421238_X1_Y1_1677466712_1677466712_0 m1_226_560# li_61_1411# PMOS_S_89421238_X1_Y1_1677466712_1677466712_0/w_0_0#
+ VSUBS PMOS_S_89421238_X1_Y1_1677466712_1677466712
XNMOS_S_25628869_X1_Y1_1677466711_1677466712_0 m1_226_560# li_61_1411# VSUBS NMOS_S_25628869_X1_Y1_1677466711_1677466712
C0 PMOS_S_89421238_X1_Y1_1677466712_1677466712_0/w_0_0# li_61_1411# 0.02fF
C1 li_61_1411# m1_226_560# 0.14fF
C2 PMOS_S_89421238_X1_Y1_1677466712_1677466712_0/w_0_0# m1_226_560# 0.55fF
C3 li_61_1411# VSUBS 0.69fF
C4 m1_226_560# VSUBS 1.33fF
C5 PMOS_S_89421238_X1_Y1_1677466712_1677466712_0/w_0_0# VSUBS 3.02fF
.ends

.subckt ANALOG_0 VN VP Y
XSTAGE2_INV_27873531_PG0_0_0_1677466713_0 m1_412_n438# m1_1088_404# VN Y VP STAGE2_INV_27873531_PG0_0_0_1677466713
XINV_21850877_PG0_0_0_1677466712_0 VN Y m1_412_n438# VP INV_21850877_PG0_0_0_1677466712
X0 VN m1_1088_404# sky130_fd_pr__cap_mim_m3_1 l=2.824e+07u w=2.897e+07u
X1 VN m1_412_n438# sky130_fd_pr__cap_mim_m3_1 l=2.824e+07u w=2.897e+07u
X2 VN Y sky130_fd_pr__cap_mim_m3_1 l=2.824e+07u w=2.897e+07u
C0 m1_412_n438# m1_1088_404# 0.21fF
C1 Y VN 5.22fF
C2 m1_412_n438# VN 8.27fF
C3 m1_412_n438# Y 2.73fF
C4 VN m1_1088_404# 4.86fF
C5 Y m1_1088_404# 2.08fF
C6 m1_1088_404# VP 12.29fF
C7 Y VP 14.86fF
C8 m1_412_n438# VP 15.87fF
C9 VN VP 12.32fF
.ends



** sch_path: /home/coold69/Documents/msvsdspwm/Week 3/xschem/analog_tb.sch
**.subckt analog_tb
X1 VN VP Y ANALOG_0
V1 VP VN 1.8
.save i(v1)
**** begin user architecture code


.lib ~/open_pdks/sources/sky130-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt
.control
save all
tran 1u 0.001
plot v(y)
.endc


.end

