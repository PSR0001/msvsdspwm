magic
tech sky130A
magscale 1 2
timestamp 1677862335
<< nwell >>
rect 0 0 1204 1512
<< pmos >>
rect 200 399 230 735
rect 286 399 316 735
rect 372 399 402 735
rect 458 399 488 735
rect 544 399 574 735
rect 630 399 660 735
rect 716 399 746 735
rect 802 399 832 735
rect 888 399 918 735
rect 974 399 1004 735
<< pdiff >>
rect 147 585 200 735
rect 147 551 155 585
rect 189 551 200 585
rect 147 517 200 551
rect 147 483 155 517
rect 189 483 200 517
rect 147 449 200 483
rect 147 415 155 449
rect 189 415 200 449
rect 147 399 200 415
rect 230 585 286 735
rect 230 551 241 585
rect 275 551 286 585
rect 230 517 286 551
rect 230 483 241 517
rect 275 483 286 517
rect 230 449 286 483
rect 230 415 241 449
rect 275 415 286 449
rect 230 399 286 415
rect 316 585 372 735
rect 316 551 327 585
rect 361 551 372 585
rect 316 517 372 551
rect 316 483 327 517
rect 361 483 372 517
rect 316 449 372 483
rect 316 415 327 449
rect 361 415 372 449
rect 316 399 372 415
rect 402 585 458 735
rect 402 551 413 585
rect 447 551 458 585
rect 402 517 458 551
rect 402 483 413 517
rect 447 483 458 517
rect 402 449 458 483
rect 402 415 413 449
rect 447 415 458 449
rect 402 399 458 415
rect 488 585 544 735
rect 488 551 499 585
rect 533 551 544 585
rect 488 517 544 551
rect 488 483 499 517
rect 533 483 544 517
rect 488 449 544 483
rect 488 415 499 449
rect 533 415 544 449
rect 488 399 544 415
rect 574 585 630 735
rect 574 551 585 585
rect 619 551 630 585
rect 574 517 630 551
rect 574 483 585 517
rect 619 483 630 517
rect 574 449 630 483
rect 574 415 585 449
rect 619 415 630 449
rect 574 399 630 415
rect 660 585 716 735
rect 660 551 671 585
rect 705 551 716 585
rect 660 517 716 551
rect 660 483 671 517
rect 705 483 716 517
rect 660 449 716 483
rect 660 415 671 449
rect 705 415 716 449
rect 660 399 716 415
rect 746 585 802 735
rect 746 551 757 585
rect 791 551 802 585
rect 746 517 802 551
rect 746 483 757 517
rect 791 483 802 517
rect 746 449 802 483
rect 746 415 757 449
rect 791 415 802 449
rect 746 399 802 415
rect 832 585 888 735
rect 832 551 843 585
rect 877 551 888 585
rect 832 517 888 551
rect 832 483 843 517
rect 877 483 888 517
rect 832 449 888 483
rect 832 415 843 449
rect 877 415 888 449
rect 832 399 888 415
rect 918 585 974 735
rect 918 551 929 585
rect 963 551 974 585
rect 918 517 974 551
rect 918 483 929 517
rect 963 483 974 517
rect 918 449 974 483
rect 918 415 929 449
rect 963 415 974 449
rect 918 399 974 415
rect 1004 585 1057 735
rect 1004 551 1015 585
rect 1049 551 1057 585
rect 1004 517 1057 551
rect 1004 483 1015 517
rect 1049 483 1057 517
rect 1004 449 1057 483
rect 1004 415 1015 449
rect 1049 415 1057 449
rect 1004 399 1057 415
<< pdiffc >>
rect 155 551 189 585
rect 155 483 189 517
rect 155 415 189 449
rect 241 551 275 585
rect 241 483 275 517
rect 241 415 275 449
rect 327 551 361 585
rect 327 483 361 517
rect 327 415 361 449
rect 413 551 447 585
rect 413 483 447 517
rect 413 415 447 449
rect 499 551 533 585
rect 499 483 533 517
rect 499 415 533 449
rect 585 551 619 585
rect 585 483 619 517
rect 585 415 619 449
rect 671 551 705 585
rect 671 483 705 517
rect 671 415 705 449
rect 757 551 791 585
rect 757 483 791 517
rect 757 415 791 449
rect 843 551 877 585
rect 843 483 877 517
rect 843 415 877 449
rect 929 551 963 585
rect 929 483 963 517
rect 929 415 963 449
rect 1015 551 1049 585
rect 1015 483 1049 517
rect 1015 415 1049 449
<< nsubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
rect 413 1361 447 1456
rect 413 1232 447 1327
rect 585 1361 619 1456
rect 585 1232 619 1327
rect 757 1361 791 1456
rect 757 1232 791 1327
rect 929 1361 963 1456
rect 929 1232 963 1327
<< nsubdiffcont >>
rect 241 1327 275 1361
rect 413 1327 447 1361
rect 585 1327 619 1361
rect 757 1327 791 1361
rect 929 1327 963 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 735 230 897
rect 286 735 316 897
rect 372 941 488 951
rect 372 907 413 941
rect 447 907 488 941
rect 372 897 488 907
rect 372 735 402 897
rect 458 735 488 897
rect 544 941 660 951
rect 544 907 585 941
rect 619 907 660 941
rect 544 897 660 907
rect 544 735 574 897
rect 630 735 660 897
rect 716 941 832 951
rect 716 907 757 941
rect 791 907 832 941
rect 716 897 832 907
rect 716 735 746 897
rect 802 735 832 897
rect 888 941 1004 951
rect 888 907 929 941
rect 963 907 1004 941
rect 888 897 1004 907
rect 888 735 918 897
rect 974 735 1004 897
rect 200 252 230 399
rect 286 252 316 399
rect 372 252 402 399
rect 458 252 488 399
rect 544 252 574 399
rect 630 252 660 399
rect 716 252 746 399
rect 802 252 832 399
rect 888 252 918 399
rect 974 252 1004 399
<< polycont >>
rect 241 907 275 941
rect 413 907 447 941
rect 585 907 619 941
rect 757 907 791 941
rect 929 907 963 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 405 1361 455 1445
rect 405 1327 413 1361
rect 447 1327 455 1361
rect 405 1243 455 1327
rect 577 1361 627 1445
rect 577 1327 585 1361
rect 619 1327 627 1361
rect 577 1243 627 1327
rect 749 1361 799 1445
rect 749 1327 757 1361
rect 791 1327 799 1361
rect 749 1243 799 1327
rect 921 1361 971 1445
rect 921 1327 929 1361
rect 963 1327 971 1361
rect 921 1243 971 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 405 941 455 1025
rect 405 907 413 941
rect 447 907 455 941
rect 405 823 455 907
rect 577 941 627 1025
rect 577 907 585 941
rect 619 907 627 941
rect 577 823 627 907
rect 749 941 799 1025
rect 749 907 757 941
rect 791 907 799 941
rect 749 823 799 907
rect 921 941 971 1025
rect 921 907 929 941
rect 963 907 971 941
rect 921 823 971 907
rect 147 585 197 773
rect 147 551 155 585
rect 189 551 197 585
rect 147 517 197 551
rect 147 483 155 517
rect 189 483 197 517
rect 147 449 197 483
rect 147 415 155 449
rect 189 415 197 449
rect 147 185 197 415
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 585 283 773
rect 233 551 241 585
rect 275 551 283 585
rect 233 517 283 551
rect 233 483 241 517
rect 275 483 283 517
rect 233 449 283 483
rect 233 415 241 449
rect 275 415 283 449
rect 233 101 283 415
rect 233 67 241 101
rect 275 67 283 101
rect 319 585 369 773
rect 319 551 327 585
rect 361 551 369 585
rect 319 517 369 551
rect 319 483 327 517
rect 361 483 369 517
rect 319 449 369 483
rect 319 415 327 449
rect 361 415 369 449
rect 319 185 369 415
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
rect 405 585 455 773
rect 405 551 413 585
rect 447 551 455 585
rect 405 517 455 551
rect 405 483 413 517
rect 447 483 455 517
rect 405 449 455 483
rect 405 415 413 449
rect 447 415 455 449
rect 405 101 455 415
rect 405 67 413 101
rect 447 67 455 101
rect 491 585 541 773
rect 491 551 499 585
rect 533 551 541 585
rect 491 517 541 551
rect 491 483 499 517
rect 533 483 541 517
rect 491 449 541 483
rect 491 415 499 449
rect 533 415 541 449
rect 491 185 541 415
rect 491 151 499 185
rect 533 151 541 185
rect 491 67 541 151
rect 577 585 627 773
rect 577 551 585 585
rect 619 551 627 585
rect 577 517 627 551
rect 577 483 585 517
rect 619 483 627 517
rect 577 449 627 483
rect 577 415 585 449
rect 619 415 627 449
rect 577 101 627 415
rect 577 67 585 101
rect 619 67 627 101
rect 663 585 713 773
rect 663 551 671 585
rect 705 551 713 585
rect 663 517 713 551
rect 663 483 671 517
rect 705 483 713 517
rect 663 449 713 483
rect 663 415 671 449
rect 705 415 713 449
rect 663 185 713 415
rect 663 151 671 185
rect 705 151 713 185
rect 663 67 713 151
rect 749 585 799 773
rect 749 551 757 585
rect 791 551 799 585
rect 749 517 799 551
rect 749 483 757 517
rect 791 483 799 517
rect 749 449 799 483
rect 749 415 757 449
rect 791 415 799 449
rect 749 101 799 415
rect 749 67 757 101
rect 791 67 799 101
rect 835 585 885 773
rect 835 551 843 585
rect 877 551 885 585
rect 835 517 885 551
rect 835 483 843 517
rect 877 483 885 517
rect 835 449 885 483
rect 835 415 843 449
rect 877 415 885 449
rect 835 185 885 415
rect 835 151 843 185
rect 877 151 885 185
rect 835 67 885 151
rect 921 585 971 773
rect 921 551 929 585
rect 963 551 971 585
rect 921 517 971 551
rect 921 483 929 517
rect 963 483 971 517
rect 921 449 971 483
rect 921 415 929 449
rect 963 415 971 449
rect 921 101 971 415
rect 921 67 929 101
rect 963 67 971 101
rect 1007 585 1057 773
rect 1007 551 1015 585
rect 1049 551 1057 585
rect 1007 517 1057 551
rect 1007 483 1015 517
rect 1049 483 1057 517
rect 1007 449 1057 483
rect 1007 415 1015 449
rect 1049 415 1057 449
rect 1007 185 1057 415
rect 1007 151 1015 185
rect 1049 151 1057 185
rect 1007 67 1057 151
<< viali >>
rect 241 1327 275 1361
rect 413 1327 447 1361
rect 585 1327 619 1361
rect 757 1327 791 1361
rect 929 1327 963 1361
rect 241 907 275 941
rect 413 907 447 941
rect 585 907 619 941
rect 757 907 791 941
rect 929 907 963 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
rect 413 67 447 101
rect 499 151 533 185
rect 585 67 619 101
rect 671 151 705 185
rect 757 67 791 101
rect 843 151 877 185
rect 929 67 963 101
rect 1015 151 1049 185
<< metal1 >>
rect 224 1370 980 1372
rect 224 1361 662 1370
rect 224 1327 241 1361
rect 275 1327 413 1361
rect 447 1327 585 1361
rect 619 1327 662 1361
rect 224 1318 662 1327
rect 714 1361 980 1370
rect 714 1327 757 1361
rect 791 1327 929 1361
rect 963 1327 980 1361
rect 714 1318 980 1327
rect 224 1316 980 1318
rect 224 941 980 952
rect 224 907 241 941
rect 275 907 413 941
rect 447 907 585 941
rect 619 907 757 941
rect 791 907 929 941
rect 963 907 980 941
rect 224 896 980 907
rect 138 194 1066 196
rect 138 185 662 194
rect 714 185 1066 194
rect 138 151 155 185
rect 189 151 327 185
rect 361 151 499 185
rect 533 151 662 185
rect 714 151 843 185
rect 877 151 1015 185
rect 1049 151 1066 185
rect 138 142 662 151
rect 714 142 1066 151
rect 138 140 1066 142
rect 224 101 980 112
rect 224 67 241 101
rect 275 67 413 101
rect 447 67 585 101
rect 619 67 757 101
rect 791 67 929 101
rect 963 67 980 101
rect 224 56 980 67
<< via1 >>
rect 662 1318 714 1370
rect 662 185 714 194
rect 662 151 671 185
rect 671 151 705 185
rect 705 151 714 185
rect 662 142 714 151
<< metal2 >>
rect 660 1370 716 1376
rect 660 1318 662 1370
rect 714 1318 716 1370
rect 660 194 716 1318
rect 660 142 662 194
rect 714 142 716 194
rect 660 136 716 142
<< end >>
