magic
tech sky130A
magscale 1 2
timestamp 1677519077
<< nwell >>
rect -18 4020 402 4202
<< locali >>
rect 491 3679 499 3713
rect 533 3679 541 3713
rect 491 3629 541 3679
rect 491 3595 499 3629
rect 533 3595 541 3629
rect 1265 3679 1273 3713
rect 1307 3679 1315 3713
rect 1265 2873 1315 3679
rect 1265 2839 1273 2873
rect 1307 2839 1315 2873
rect 1093 2201 1143 2688
rect 1093 2167 1101 2201
rect 1135 2167 1143 2201
<< viali >>
rect 499 3679 533 3713
rect 499 3595 533 3629
rect 1273 3679 1307 3713
rect 1273 2839 1307 2873
rect 1101 2167 1135 2201
<< metal1 >>
rect -18 4020 402 4202
rect 430 3713 550 3724
rect 430 3679 499 3713
rect 533 3679 550 3713
rect 430 3668 550 3679
rect 1256 3713 1462 3724
rect 1256 3679 1273 3713
rect 1307 3679 1462 3713
rect 1256 3668 1462 3679
rect 482 3638 1494 3640
rect 482 3629 1436 3638
rect 482 3595 499 3629
rect 533 3595 1436 3629
rect 482 3586 1436 3595
rect 1488 3586 1494 3638
rect 482 3584 1494 3586
rect 484 3050 1408 3052
rect 484 2998 490 3050
rect 542 2998 834 3050
rect 886 2998 1350 3050
rect 1402 2998 1408 3050
rect 484 2996 1408 2998
rect 226 2882 290 2884
rect 226 2830 232 2882
rect 284 2830 290 2882
rect 226 2828 290 2830
rect 1118 2873 1324 2884
rect 1118 2839 1273 2873
rect 1307 2839 1324 2873
rect 1118 2828 1324 2839
rect 1430 2882 1494 2884
rect 1430 2830 1436 2882
rect 1488 2830 1494 2882
rect 1430 2828 1494 2830
rect 1084 2210 1322 2212
rect 1084 2201 1264 2210
rect 1084 2167 1101 2201
rect 1135 2167 1264 2201
rect 1084 2158 1264 2167
rect 1316 2158 1322 2210
rect 1084 2156 1322 2158
rect 656 1874 946 1876
rect 656 1822 662 1874
rect 714 1822 946 1874
rect 656 1820 946 1822
rect 430 1454 720 1456
rect 430 1402 662 1454
rect 714 1402 720 1454
rect 430 1400 720 1402
rect 914 1370 1290 1372
rect 914 1318 920 1370
rect 972 1318 1290 1370
rect 914 1316 1290 1318
rect 1430 1370 1494 1372
rect 1430 1318 1436 1370
rect 1488 1318 1494 1370
rect 1430 1316 1494 1318
rect 430 614 548 616
rect 430 562 490 614
rect 542 562 548 614
rect 430 560 548 562
<< via1 >>
rect 1436 3586 1488 3638
rect 490 2998 542 3050
rect 834 2998 886 3050
rect 1350 2998 1402 3050
rect 232 2830 284 2882
rect 1436 2830 1488 2882
rect 1264 2158 1316 2210
rect 662 1822 714 1874
rect 662 1402 714 1454
rect 920 1318 972 1370
rect 1436 1318 1488 1370
rect 490 562 542 614
<< metal2 >>
rect 1434 3638 1490 3644
rect 1434 3586 1436 3638
rect 1488 3586 1490 3638
rect 488 3050 544 3056
rect 488 2998 490 3050
rect 542 2998 544 3050
rect 488 2992 544 2998
rect 832 3050 888 3056
rect 832 2998 834 3050
rect 886 2998 888 3050
rect 832 2992 888 2998
rect 1348 3050 1404 3056
rect 1348 2998 1350 3050
rect 1402 2998 1404 3050
rect 1348 2992 1404 2998
rect 230 2882 286 2888
rect 230 2830 232 2882
rect 284 2830 286 2882
rect 230 2548 286 2830
rect 1434 2882 1490 3586
rect 1434 2830 1436 2882
rect 1488 2830 1490 2882
rect 230 2483 286 2492
rect 918 2548 974 2557
rect 918 2483 974 2492
rect 1262 2210 1318 2216
rect 1262 2158 1264 2210
rect 1316 2158 1318 2210
rect 660 1874 716 1880
rect 660 1822 662 1874
rect 714 1822 716 1874
rect 144 1792 200 1801
rect 144 1344 200 1736
rect 660 1454 716 1822
rect 832 1792 888 1801
rect 832 1727 888 1736
rect 660 1402 662 1454
rect 714 1402 716 1454
rect 660 1396 716 1402
rect 918 1370 974 1376
rect 918 1318 920 1370
rect 972 1318 974 1370
rect 488 1036 544 1045
rect 488 614 544 980
rect 918 1036 974 1318
rect 918 971 974 980
rect 1262 1036 1318 2158
rect 1434 1370 1490 2830
rect 1520 1792 1576 1801
rect 1520 1727 1576 1736
rect 1434 1318 1436 1370
rect 1488 1318 1490 1370
rect 1434 1312 1490 1318
rect 1262 971 1318 980
rect 488 562 490 614
rect 542 562 544 614
rect 488 556 544 562
rect 144 280 200 289
rect 144 215 200 224
<< via2 >>
rect 230 2492 286 2548
rect 918 2492 974 2548
rect 144 1736 200 1792
rect 832 1736 888 1792
rect 488 980 544 1036
rect 918 980 974 1036
rect 1520 1736 1576 1792
rect 1262 980 1318 1036
rect 144 224 200 280
<< metal3 >>
rect 225 2548 291 2600
rect 225 2492 230 2548
rect 286 2492 291 2548
rect 225 2440 291 2492
rect 602 2548 979 2600
rect 602 2492 918 2548
rect 974 2492 979 2548
rect 602 2440 979 2492
rect 139 1792 258 1844
rect 139 1736 144 1792
rect 200 1736 258 1792
rect 139 1684 258 1736
rect 602 1792 1581 1844
rect 602 1736 832 1792
rect 888 1736 1520 1792
rect 1576 1736 1581 1792
rect 602 1684 1581 1736
rect 483 1036 592 1088
rect 483 980 488 1036
rect 544 980 592 1036
rect 483 928 592 980
rect 913 1036 979 1088
rect 913 980 918 1036
rect 974 980 979 1036
rect 913 928 979 980
rect 1257 1036 1323 1088
rect 1257 980 1262 1036
rect 1318 980 1323 1036
rect 1257 928 1323 980
rect 139 280 592 332
rect 139 224 144 280
rect 200 224 592 280
rect 139 172 592 224
rect 946 172 1184 332
use CAP_2T_9576091_1677407591  CAP_2T_9576091_1677407591_0
timestamp 1677423745
transform 1 0 1118 0 1 0
box 53 166 463 1088
use CAP_2T_9576091_1677407591  CAP_2T_9576091_1677407591_1
timestamp 1677423745
transform -1 0 688 0 1 1512
box 53 166 463 1088
use CAP_2T_9576091_1677407591  CAP_2T_9576091_1677407591_2
timestamp 1677423745
transform 1 0 516 0 1 0
box 53 166 463 1088
use INV_21850877_0_0_1677407590  INV_21850877_0_0_1677407590_0
timestamp 1677423745
transform 1 0 688 0 1 1260
box 0 30 516 3024
use NMOS_S_25628869_X1_Y1_1677407592  NMOS_S_25628869_X1_Y1_1677407592_0
timestamp 1677423745
transform -1 0 516 0 -1 1512
box 52 56 395 1482
use NMOS_S_25628869_X1_Y1_1677407592  NMOS_S_25628869_X1_Y1_1677407592_1
timestamp 1677423745
transform 1 0 1204 0 1 1260
box 52 56 395 1482
use PMOS_S_89421238_X1_Y1_1677407593  PMOS_S_89421238_X1_Y1_1677407593_0
timestamp 1677423745
transform -1 0 1720 0 1 2772
box 0 0 516 1512
use PMOS_S_89421238_X1_Y1_1677407593  PMOS_S_89421238_X1_Y1_1677407593_1
timestamp 1677423745
transform 1 0 172 0 1 2772
box 0 0 516 1512
<< labels >>
rlabel space 636 250 636 250 1 VN
port 1 n
rlabel metal1 1194 2176 1194 2176 1 Y
port 3 n
<< end >>
