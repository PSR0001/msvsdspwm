magic
tech sky130A
magscale 1 2
timestamp 1676537953
<< nwell >>
rect -208 2020 3398 2704
rect -208 1946 542 2020
rect 574 1946 3398 2020
rect -208 1792 3398 1946
<< metal1 >>
rect -210 2710 3396 2858
rect -202 2306 -80 2710
rect 956 2554 2256 2646
rect 66 2420 152 2424
rect 66 2362 82 2420
rect 138 2362 152 2420
rect 66 2358 152 2362
rect 666 2420 752 2424
rect 666 2362 680 2420
rect 736 2362 752 2420
rect 666 2358 752 2362
rect 958 2306 1068 2554
rect 1868 2422 1954 2426
rect 1268 2416 1354 2422
rect 1268 2358 1284 2416
rect 1340 2358 1354 2416
rect 1868 2364 1884 2422
rect 1940 2364 1954 2422
rect 1868 2360 1954 2364
rect 1268 2356 1354 2358
rect 2146 2308 2256 2554
rect 2468 2418 2554 2422
rect 2468 2360 2482 2418
rect 2538 2360 2554 2418
rect 2468 2356 2554 2360
rect 3066 2420 3152 2424
rect 3066 2362 3084 2420
rect 3140 2362 3152 2420
rect 3066 2358 3152 2362
rect 3312 2310 3388 2710
rect -202 2128 82 2306
rect 136 2130 686 2306
rect 738 2130 1288 2306
rect 1340 2130 1890 2306
rect 1942 2132 2492 2308
rect 2538 2132 3088 2308
rect 3138 2132 3388 2310
rect -202 2126 -80 2128
rect 66 2074 152 2080
rect 66 2016 82 2074
rect 138 2016 152 2074
rect 66 2014 152 2016
rect 668 2074 754 2078
rect 668 2016 682 2074
rect 738 2016 754 2074
rect 668 2012 754 2016
rect 1268 2074 1354 2078
rect 1268 2016 1282 2074
rect 1338 2016 1354 2074
rect 1268 2012 1354 2016
rect 1560 1722 1666 2130
rect 1868 2074 1954 2080
rect 1868 2016 1884 2074
rect 1940 2016 1954 2074
rect 1868 2014 1954 2016
rect 2470 2076 2556 2080
rect 2470 2018 2484 2076
rect 2540 2018 2556 2076
rect 2470 2014 2556 2018
rect 3068 2078 3154 2082
rect 3068 2020 3082 2078
rect 3138 2020 3154 2078
rect 3068 2016 3154 2020
rect -184 1644 3406 1722
rect -180 1396 -110 1644
rect 66 1502 152 1504
rect 66 1444 82 1502
rect 138 1444 152 1502
rect 66 1438 152 1444
rect 664 1500 750 1504
rect 664 1442 678 1500
rect 734 1442 750 1500
rect 664 1438 750 1442
rect 960 1396 1042 1644
rect 1264 1504 1350 1506
rect 1264 1446 1278 1504
rect 1334 1446 1350 1504
rect 1264 1440 1350 1446
rect 1868 1498 1954 1502
rect 1868 1440 1886 1498
rect 1942 1440 1954 1498
rect 1868 1436 1954 1440
rect 2470 1498 2556 1502
rect 2470 1440 2484 1498
rect 2540 1440 2556 1498
rect 3068 1500 3154 1508
rect 3068 1442 3082 1500
rect 3138 1442 3154 1500
rect 2470 1436 2556 1440
rect -180 1220 84 1396
rect 136 1360 682 1396
rect 136 1286 350 1360
rect 424 1286 682 1360
rect 136 1220 682 1286
rect 736 1220 1282 1396
rect 1334 1224 1886 1396
rect 1940 1222 2486 1396
rect 2540 1354 3084 1400
rect 2540 1280 2774 1354
rect 2848 1280 3084 1354
rect 1262 1178 1348 1182
rect 66 1172 152 1178
rect 66 1114 82 1172
rect 138 1114 152 1172
rect 66 1112 152 1114
rect 664 1174 750 1178
rect 664 1116 680 1174
rect 736 1116 750 1174
rect 1262 1120 1276 1178
rect 1332 1120 1348 1178
rect 1262 1116 1348 1120
rect 1870 1174 1956 1178
rect 1870 1116 1884 1174
rect 1940 1116 1956 1174
rect 664 1112 750 1116
rect 1870 1112 1956 1116
rect 2160 970 2246 1222
rect 2540 1220 3084 1280
rect 3138 1224 3306 1400
rect 3066 1180 3152 1182
rect 2472 1174 2558 1178
rect 2472 1116 2482 1174
rect 2538 1116 2558 1174
rect 3066 1122 3086 1180
rect 3142 1122 3152 1180
rect 3066 1116 3152 1122
rect 2472 1112 2558 1116
rect 3216 970 3302 1224
rect -206 794 3400 970
<< via1 >>
rect 82 2362 138 2420
rect 680 2362 736 2420
rect 1284 2358 1340 2416
rect 1884 2364 1940 2422
rect 2482 2360 2538 2418
rect 3084 2362 3140 2420
rect 82 2016 138 2074
rect 682 2016 738 2074
rect 1282 2016 1338 2074
rect 1884 2016 1940 2074
rect 2484 2018 2540 2076
rect 3082 2020 3138 2078
rect 82 1444 138 1502
rect 678 1442 734 1500
rect 1278 1446 1334 1504
rect 1886 1440 1942 1498
rect 2484 1440 2540 1498
rect 3082 1442 3138 1500
rect 350 1286 424 1360
rect 2774 1280 2848 1354
rect 82 1114 138 1172
rect 680 1116 736 1174
rect 1276 1120 1332 1178
rect 1884 1116 1940 1174
rect 2482 1116 2538 1174
rect 3086 1122 3142 1180
<< metal2 >>
rect 66 2420 152 2424
rect 66 2362 82 2420
rect 138 2362 152 2420
rect 66 2358 152 2362
rect 666 2420 752 2424
rect 1868 2422 1954 2426
rect 666 2362 680 2420
rect 736 2362 752 2420
rect 666 2358 752 2362
rect 1268 2416 1354 2422
rect 1268 2358 1284 2416
rect 1340 2358 1354 2416
rect 1868 2364 1884 2422
rect 1940 2364 1954 2422
rect 1868 2360 1954 2364
rect 2468 2418 2554 2422
rect 2468 2360 2482 2418
rect 2538 2360 2554 2418
rect 90 2080 128 2358
rect 66 2074 152 2080
rect 690 2078 728 2358
rect 1268 2356 1354 2358
rect 1290 2078 1328 2356
rect 1894 2080 1932 2360
rect 2468 2356 2554 2360
rect 3066 2420 3152 2424
rect 3066 2362 3084 2420
rect 3140 2362 3152 2420
rect 3066 2358 3152 2362
rect 2494 2080 2532 2356
rect 3094 2082 3132 2358
rect 66 2016 82 2074
rect 138 2016 152 2074
rect 66 2014 152 2016
rect 668 2074 754 2078
rect 668 2016 682 2074
rect 738 2016 754 2074
rect 90 1504 128 2014
rect 668 2012 754 2016
rect 1268 2074 1354 2078
rect 1268 2016 1282 2074
rect 1338 2016 1354 2074
rect 1268 2012 1354 2016
rect 1868 2074 1954 2080
rect 1868 2016 1884 2074
rect 1940 2016 1954 2074
rect 1868 2014 1954 2016
rect 2470 2076 2556 2080
rect 2470 2018 2484 2076
rect 2540 2018 2556 2076
rect 2470 2014 2556 2018
rect 3068 2078 3154 2082
rect 3068 2020 3082 2078
rect 3138 2020 3154 2078
rect 3068 2016 3154 2020
rect 690 1504 728 2012
rect 1290 1506 1328 2012
rect 1264 1504 1350 1506
rect 66 1502 152 1504
rect 66 1444 82 1502
rect 138 1444 152 1502
rect 66 1438 152 1444
rect 664 1500 750 1504
rect 664 1442 678 1500
rect 734 1442 750 1500
rect 664 1438 750 1442
rect 1264 1446 1278 1504
rect 1334 1446 1350 1504
rect 1894 1502 1932 2014
rect 2494 1502 2532 2014
rect 3094 1508 3132 2016
rect 1264 1440 1350 1446
rect 1868 1498 1954 1502
rect 1868 1440 1886 1498
rect 1942 1440 1954 1498
rect 90 1178 128 1438
rect 344 1360 432 1368
rect 344 1286 350 1360
rect 424 1286 432 1360
rect 66 1172 152 1178
rect 66 1114 82 1172
rect 138 1114 152 1172
rect 66 1112 152 1114
rect 344 1064 432 1286
rect 690 1178 728 1438
rect 1290 1182 1328 1440
rect 1868 1436 1954 1440
rect 2470 1498 2556 1502
rect 2470 1440 2484 1498
rect 2540 1440 2556 1498
rect 3068 1500 3154 1508
rect 3068 1442 3082 1500
rect 3138 1442 3154 1500
rect 2470 1436 2556 1440
rect 1262 1178 1348 1182
rect 1894 1178 1932 1436
rect 2494 1178 2532 1436
rect 2768 1354 2856 1366
rect 2768 1280 2774 1354
rect 2848 1280 2856 1354
rect 664 1174 750 1178
rect 664 1116 680 1174
rect 736 1116 750 1174
rect 1262 1120 1276 1178
rect 1332 1120 1348 1178
rect 1262 1116 1348 1120
rect 1870 1174 1956 1178
rect 1870 1116 1884 1174
rect 1940 1116 1956 1174
rect 664 1112 750 1116
rect 1870 1112 1956 1116
rect 2472 1174 2558 1178
rect 2472 1116 2482 1174
rect 2538 1116 2558 1174
rect 2472 1112 2558 1116
rect 2768 1064 2856 1280
rect 3094 1182 3132 1442
rect 3066 1180 3152 1182
rect 3066 1122 3086 1180
rect 3142 1122 3152 1180
rect 3066 1116 3152 1122
rect 344 980 2856 1064
use sky130_fd_pr__nfet_01v8_648S5X  XM1
timestamp 1676522790
transform 1 0 109 0 1 1308
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM2
timestamp 1676522790
transform 1 0 709 0 1 1308
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM3
timestamp 1676522790
transform 1 0 1307 0 1 1312
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM4
timestamp 1676522790
transform 1 0 1913 0 1 1308
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM5
timestamp 1676522790
transform 1 0 3111 0 1 1312
box -211 -310 211 310
use sky130_fd_pr__nfet_01v8_648S5X  XM6
timestamp 1676522790
transform 1 0 2513 0 1 1308
box -211 -310 211 310
use sky130_fd_pr__pfet_01v8_XGS3BL  XM7
timestamp 1676403207
transform 1 0 1311 0 1 2217
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM8
timestamp 1676403207
transform 1 0 1913 0 1 2221
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM9
timestamp 1676403207
transform 1 0 109 0 1 2219
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM10
timestamp 1676403207
transform 1 0 711 0 1 2219
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM11
timestamp 1676403207
transform 1 0 3111 0 1 2221
box -211 -319 211 319
use sky130_fd_pr__pfet_01v8_XGS3BL  XM12
timestamp 1676403207
transform 1 0 2511 0 1 2219
box -211 -319 211 319
<< labels >>
flabel metal1 1286 860 1286 860 0 FreeSans 640 0 0 0 GND
port 9 nsew
flabel metal1 1446 2772 1446 2772 0 FreeSans 640 0 0 0 VDD
port 8 nsew
rlabel metal2 112 1756 112 1756 1 A
port 1 n
rlabel metal2 706 1754 706 1754 1 C
port 2 n
rlabel metal2 1308 1748 1308 1748 1 E
port 3 n
rlabel metal2 1912 1752 1912 1752 1 F
port 4 n
rlabel metal2 2514 1754 2514 1754 1 D
port 5 n
rlabel metal2 3110 1758 3110 1758 1 B
port 6 n
rlabel metal1 3370 1684 3370 1684 1 Y
port 7 n
<< end >>
