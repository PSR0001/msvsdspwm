magic
tech sky130A
magscale 1 2
timestamp 1678383033
<< locali >>
rect 577 2419 585 2453
rect 619 2419 627 2453
rect 61 1579 69 1613
rect 103 1579 111 1613
rect 61 1445 111 1579
rect 61 1411 69 1445
rect 103 1411 111 1445
rect 577 1445 627 2419
rect 577 1411 585 1445
rect 619 1411 627 1445
rect 921 1579 929 1613
rect 963 1579 971 1613
rect 921 1445 971 1579
rect 921 1411 929 1445
rect 963 1411 971 1445
rect 577 605 627 1411
rect 577 571 585 605
rect 619 571 627 605
<< viali >>
rect 585 2419 619 2453
rect 69 1579 103 1613
rect 69 1411 103 1445
rect 585 1411 619 1445
rect 929 1579 963 1613
rect 929 1411 963 1445
rect 585 571 619 605
<< metal1 >>
rect 258 2453 636 2464
rect 258 2419 585 2453
rect 619 2419 636 2453
rect 258 2408 636 2419
rect 742 2462 806 2464
rect 742 2410 748 2462
rect 800 2410 806 2462
rect 742 2408 806 2410
rect 312 1790 720 1792
rect 312 1738 318 1790
rect 370 1738 662 1790
rect 714 1738 720 1790
rect 312 1736 720 1738
rect 52 1613 120 1624
rect 52 1579 69 1613
rect 103 1579 120 1613
rect 52 1568 120 1579
rect 912 1613 980 1624
rect 912 1579 929 1613
rect 963 1579 980 1613
rect 912 1568 980 1579
rect 52 1445 120 1456
rect 52 1411 69 1445
rect 103 1411 120 1445
rect 52 1400 120 1411
rect 568 1445 774 1456
rect 568 1411 585 1445
rect 619 1411 774 1445
rect 568 1400 774 1411
rect 912 1445 980 1456
rect 912 1411 929 1445
rect 963 1411 980 1445
rect 912 1400 980 1411
rect 258 605 636 616
rect 258 571 585 605
rect 619 571 636 605
rect 258 560 636 571
rect 742 614 806 616
rect 742 562 748 614
rect 800 562 806 614
rect 742 560 806 562
rect 312 278 720 280
rect 312 226 318 278
rect 370 226 662 278
rect 714 226 720 278
rect 312 224 720 226
<< via1 >>
rect 748 2410 800 2462
rect 318 1738 370 1790
rect 662 1738 714 1790
rect 748 562 800 614
rect 318 226 370 278
rect 662 226 714 278
<< metal2 >>
rect 746 2462 802 2468
rect 746 2410 748 2462
rect 800 2410 802 2462
rect 316 1790 372 1796
rect 316 1738 318 1790
rect 370 1738 372 1790
rect 316 1732 372 1738
rect 660 1790 716 1796
rect 660 1738 662 1790
rect 714 1738 716 1790
rect 660 1732 716 1738
rect 746 614 802 2410
rect 746 562 748 614
rect 800 562 802 614
rect 746 556 802 562
rect 316 278 372 284
rect 316 226 318 278
rect 370 226 372 278
rect 316 220 372 226
rect 660 278 716 284
rect 660 226 662 278
rect 714 226 716 278
rect 660 220 716 226
use NMOS_S_94657632_X1_Y1_1678381962_1678381963  NMOS_S_94657632_X1_Y1_1678381962_1678381963_0
timestamp 1678383033
transform 1 0 0 0 -1 1512
box 52 56 395 1482
use NMOS_S_94657632_X1_Y1_1678381962_1678381963  NMOS_S_94657632_X1_Y1_1678381962_1678381963_1
timestamp 1678383033
transform -1 0 1032 0 -1 1512
box 52 56 395 1482
use PMOS_S_13339638_X1_Y1_1678381963_1678381963  PMOS_S_13339638_X1_Y1_1678381963_1678381963_0
timestamp 1678383033
transform 1 0 0 0 1 1512
box 0 0 516 1512
use PMOS_S_13339638_X1_Y1_1678381963_1678381963  PMOS_S_13339638_X1_Y1_1678381963_1678381963_1
timestamp 1678383033
transform -1 0 1032 0 1 1512
box 0 0 516 1512
<< end >>
