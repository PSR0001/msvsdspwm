magic
tech sky130A
magscale 1 2
timestamp 1677862335
<< metal1 >>
rect 484 1790 720 1792
rect 484 1738 490 1790
rect 542 1738 662 1790
rect 714 1738 720 1790
rect 484 1736 720 1738
rect 1602 1790 1752 1792
rect 1602 1738 1608 1790
rect 1660 1738 1694 1790
rect 1746 1738 1752 1790
rect 1602 1736 1752 1738
rect 2806 1790 2956 1792
rect 2806 1738 2812 1790
rect 2864 1738 2898 1790
rect 2950 1738 2956 1790
rect 2806 1736 2956 1738
rect 1258 1538 1580 1540
rect 1258 1486 1264 1538
rect 1316 1486 1522 1538
rect 1574 1486 1580 1538
rect 1258 1484 1580 1486
rect 946 1454 1322 1456
rect 946 1402 1264 1454
rect 1316 1402 1322 1454
rect 946 1400 1322 1402
rect 570 1286 720 1288
rect 570 1234 576 1286
rect 628 1234 662 1286
rect 714 1234 720 1286
rect 570 1232 720 1234
<< via1 >>
rect 490 1738 542 1790
rect 662 1738 714 1790
rect 1608 1738 1660 1790
rect 1694 1738 1746 1790
rect 2812 1738 2864 1790
rect 2898 1738 2950 1790
rect 1264 1486 1316 1538
rect 1522 1486 1574 1538
rect 1264 1402 1316 1454
rect 576 1234 628 1286
rect 662 1234 714 1286
<< metal2 >>
rect 488 1790 544 1796
rect 488 1738 490 1790
rect 542 1738 544 1790
rect 316 1540 372 1549
rect 316 1475 372 1484
rect 488 28 544 1738
rect 574 1792 630 1801
rect 574 1286 630 1736
rect 660 1790 716 1796
rect 660 1738 662 1790
rect 714 1738 716 1790
rect 660 1732 716 1738
rect 1606 1790 1662 1796
rect 1606 1738 1608 1790
rect 1660 1738 1662 1790
rect 1262 1538 1318 1544
rect 1262 1486 1264 1538
rect 1316 1486 1318 1538
rect 1262 1454 1318 1486
rect 1520 1538 1576 1544
rect 1520 1486 1522 1538
rect 1574 1486 1576 1538
rect 1520 1480 1576 1486
rect 1262 1402 1264 1454
rect 1316 1402 1318 1454
rect 1262 1396 1318 1402
rect 574 1234 576 1286
rect 628 1234 630 1286
rect 574 1228 630 1234
rect 660 1286 716 1292
rect 660 1234 662 1286
rect 714 1234 716 1286
rect 660 1228 716 1234
rect 488 -37 544 -28
rect 1606 28 1662 1738
rect 1692 1790 1748 1796
rect 1692 1738 1694 1790
rect 1746 1738 1748 1790
rect 1692 1732 1748 1738
rect 2810 1790 2866 1796
rect 2810 1738 2812 1790
rect 2864 1738 2866 1790
rect 2638 1540 2694 1549
rect 2638 1475 2694 1484
rect 1692 1288 1748 1297
rect 1692 1223 1748 1232
rect 1606 -37 1662 -28
rect 2810 28 2866 1738
rect 2896 1790 2952 1796
rect 2896 1738 2898 1790
rect 2950 1738 2952 1790
rect 2896 1732 2952 1738
rect 2896 1288 2952 1297
rect 2896 1223 2952 1232
rect 2810 -37 2866 -28
<< via2 >>
rect 316 1484 372 1540
rect 574 1736 630 1792
rect 488 -28 544 28
rect 2638 1484 2694 1540
rect 1692 1232 1748 1288
rect 1606 -28 1662 28
rect 2896 1232 2952 1288
rect 2810 -28 2866 28
<< metal3 >>
rect -80 1796 3520 1844
rect -80 1792 1744 1796
rect -80 1736 574 1792
rect 630 1736 1744 1792
rect -80 1732 1744 1736
rect 1808 1732 2336 1796
rect 2400 1732 2928 1796
rect 2992 1732 3520 1796
rect -80 1684 3520 1732
rect 311 1540 2699 1592
rect 311 1484 316 1540
rect 372 1484 2638 1540
rect 2694 1484 2699 1540
rect 311 1432 2699 1484
rect 1687 1292 1809 1340
rect 1687 1288 1744 1292
rect 1687 1232 1692 1288
rect 1687 1228 1744 1232
rect 1808 1228 1809 1292
rect 1687 1180 1809 1228
rect 2891 1292 2993 1340
rect 2891 1288 2928 1292
rect 2891 1232 2896 1288
rect 2891 1228 2928 1232
rect 2992 1228 2993 1292
rect 2891 1180 2993 1228
rect -80 32 3520 80
rect -80 -32 -32 32
rect 32 28 3520 32
rect 32 -28 488 28
rect 544 -28 1606 28
rect 1662 -28 2810 28
rect 2866 -28 3520 28
rect 32 -32 3520 -28
rect -80 -80 3520 -32
<< via3 >>
rect 1744 1732 1808 1796
rect 2336 1732 2400 1796
rect 2928 1732 2992 1796
rect 1744 1288 1808 1292
rect 1744 1232 1748 1288
rect 1748 1232 1808 1288
rect 1744 1228 1808 1232
rect 2928 1288 2992 1292
rect 2928 1232 2952 1288
rect 2952 1232 2992 1288
rect 2928 1228 2992 1232
rect -32 -32 32 32
<< metal4 >>
rect -118 32 118 1882
rect 1658 1796 1894 1797
rect 1658 1732 1744 1796
rect 1808 1732 1894 1796
rect 1658 1292 1894 1732
rect 1658 1228 1744 1292
rect 1808 1228 1894 1292
rect 1658 1227 1894 1228
rect 2250 1796 2486 1882
rect 2250 1732 2336 1796
rect 2400 1732 2486 1796
rect -118 -32 -32 32
rect 32 -32 118 32
rect -118 -118 118 -32
rect 2250 -118 2486 1732
rect 2842 1796 3078 1797
rect 2842 1732 2928 1796
rect 2992 1732 3078 1796
rect 2842 1292 3078 1732
rect 2842 1228 2928 1292
rect 2992 1228 3078 1292
rect 2842 1227 3078 1228
use INV_8026114_PG0_0_0_1677862246  INV_8026114_PG0_0_0_1677862246_0
timestamp 1677862335
transform 1 0 0 0 1 0
box 0 30 1204 3024
use STAGE2_INV_31651850_PG0_0_0_1677862247  STAGE2_INV_31651850_PG0_0_0_1677862247_0
timestamp 1677862335
transform -1 0 3612 0 1 0
box 0 30 2408 3024
<< labels >>
flabel metal1 s 602 1428 602 1428 0 FreeSerif 0 0 0 0 Y
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal3 s 1748 1260 1748 1260 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 VN
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
flabel metal1 s 1677 1764 1677 1764 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VP
<< end >>
