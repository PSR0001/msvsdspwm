magic
tech sky130A
magscale 1 2
timestamp 1677862335
<< locali >>
rect 1093 2419 1101 2453
rect 1135 2419 1143 2453
rect 1093 1445 1143 2419
rect 1093 1411 1101 1445
rect 1135 1411 1143 1445
rect 1093 605 1143 1411
rect 1093 571 1101 605
rect 1135 571 1143 605
<< viali >>
rect 1101 2419 1135 2453
rect 1101 1411 1135 1445
rect 1101 571 1135 605
<< metal1 >>
rect 946 2453 1152 2464
rect 946 2419 1101 2453
rect 1135 2419 1152 2453
rect 946 2408 1152 2419
rect 2032 2462 2096 2464
rect 2032 2410 2038 2462
rect 2090 2410 2096 2462
rect 2032 2408 2096 2410
rect 914 1622 978 1624
rect 914 1570 920 1622
rect 972 1570 978 1622
rect 914 1568 978 1570
rect 2118 1622 2182 1624
rect 2118 1570 2124 1622
rect 2176 1570 2182 1622
rect 2118 1568 2182 1570
rect 914 1454 978 1456
rect 914 1402 920 1454
rect 972 1402 978 1454
rect 914 1400 978 1402
rect 1084 1445 1462 1456
rect 1084 1411 1101 1445
rect 1135 1411 1462 1445
rect 1084 1400 1462 1411
rect 2118 1454 2182 1456
rect 2118 1402 2124 1454
rect 2176 1402 2182 1454
rect 2118 1400 2182 1402
rect 946 605 1152 616
rect 946 571 1101 605
rect 1135 571 1152 605
rect 946 560 1152 571
rect 2032 614 2096 616
rect 2032 562 2038 614
rect 2090 562 2096 614
rect 2032 560 2096 562
<< via1 >>
rect 2038 2410 2090 2462
rect 920 1570 972 1622
rect 2124 1570 2176 1622
rect 920 1402 972 1454
rect 2124 1402 2176 1454
rect 2038 562 2090 614
<< metal2 >>
rect 2036 2462 2092 2468
rect 2036 2410 2038 2462
rect 2090 2410 2092 2462
rect 918 1622 974 1628
rect 918 1570 920 1622
rect 972 1570 974 1622
rect 918 1454 974 1570
rect 918 1402 920 1454
rect 972 1402 974 1454
rect 918 1396 974 1402
rect 2036 614 2092 2410
rect 2122 1622 2178 1628
rect 2122 1570 2124 1622
rect 2176 1570 2178 1622
rect 2122 1454 2178 1570
rect 2122 1402 2124 1454
rect 2176 1402 2178 1454
rect 2122 1396 2178 1402
rect 2036 562 2038 614
rect 2090 562 2092 614
rect 2036 556 2092 562
use NMOS_S_4459928_X5_Y1_1677862245_1677862247  NMOS_S_4459928_X5_Y1_1677862245_1677862247_0
timestamp 1677862335
transform 1 0 0 0 -1 1512
box 121 56 1083 1482
use NMOS_S_4459928_X5_Y1_1677862245_1677862247  NMOS_S_4459928_X5_Y1_1677862245_1677862247_1
timestamp 1677862335
transform 1 0 1204 0 -1 1512
box 121 56 1083 1482
use PMOS_S_62253992_X5_Y1_1677862246_1677862247  PMOS_S_62253992_X5_Y1_1677862246_1677862247_0
timestamp 1677862335
transform 1 0 0 0 1 1512
box 0 0 1204 1512
use PMOS_S_62253992_X5_Y1_1677862246_1677862247  PMOS_S_62253992_X5_Y1_1677862246_1677862247_1
timestamp 1677862335
transform 1 0 1204 0 1 1512
box 0 0 1204 1512
<< end >>
