X1 in out net1 GND inverter
V1 net1 GND 1.8
.save i(v1)
V2 in GND pulse(0 1.8 1n 1n 1n 4n 10n)
.save i(v2)
**** begin user architecture code

.lib ~/open_pdks/sources/sky130-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt
.control
save all
tran 1n 20n
plot v(in) v(out)
.endc

.subckt INV vin vout vdd vss
XM2 vout vin vss vss sky130_fd_pr__nfet_01v8 L=0.15 W=4.2 nf=2 
XM3 vout vin vdd vdd sky130_fd_pr__pfet_01v8 L=0.15 W=8.4 nf=2
.ends
.GLOBAL GND
.end
