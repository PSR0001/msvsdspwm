magic
tech sky130A
magscale 1 2
timestamp 1678376823
<< error_s >>
rect 2004 1568 2012 1624
rect 2032 1568 2040 1624
rect 2520 1568 2528 1624
rect 2548 1568 2556 1624
rect 2520 1400 2528 1456
rect 2548 1400 2556 1456
<< nwell >>
rect 1016 1508 1458 1790
<< locali >>
rect 1265 1747 1273 1781
rect 1307 1747 1315 1781
rect 491 1579 499 1613
rect 533 1579 541 1613
rect 491 1529 541 1579
rect 491 1495 499 1529
rect 533 1495 541 1529
rect 1179 1327 1187 1361
rect 1221 1327 1229 1361
rect 1179 1277 1229 1327
rect 1179 1243 1187 1277
rect 1221 1243 1229 1277
rect 1265 17 1315 1747
rect 2641 1579 2649 1613
rect 2683 1579 2691 1613
rect 2125 1495 2133 1529
rect 2167 1495 2175 1529
rect 2125 1445 2175 1495
rect 2125 1411 2133 1445
rect 2167 1411 2175 1445
rect 1265 -17 1273 17
rect 1307 -17 1315 17
rect 2641 17 2691 1579
rect 2641 -17 2649 17
rect 2683 -17 2691 17
<< viali >>
rect 1273 1747 1307 1781
rect 499 1579 533 1613
rect 499 1495 533 1529
rect 1187 1327 1221 1361
rect 1187 1243 1221 1277
rect 2649 1579 2683 1613
rect 2133 1495 2167 1529
rect 2133 1411 2167 1445
rect 1273 -17 1307 17
rect 2649 -17 2683 17
<< metal1 >>
rect 312 2882 376 2884
rect 312 2830 318 2882
rect 370 2830 376 2882
rect 312 2828 376 2830
rect 828 2882 892 2884
rect 828 2830 834 2882
rect 886 2830 892 2882
rect 828 2828 892 2830
rect 474 2428 552 2486
rect 1010 2448 1066 2494
rect 1256 1790 1408 1792
rect 1256 1781 1350 1790
rect 1256 1747 1273 1781
rect 1307 1747 1350 1781
rect 1256 1738 1350 1747
rect 1402 1738 1408 1790
rect 1256 1736 1408 1738
rect 226 1706 290 1708
rect 226 1654 232 1706
rect 284 1654 290 1706
rect 226 1652 290 1654
rect 430 1652 774 1708
rect 482 1613 550 1624
rect 482 1579 499 1613
rect 533 1579 550 1613
rect 482 1568 550 1579
rect 828 1622 892 1624
rect 828 1570 834 1622
rect 886 1570 892 1622
rect 828 1568 892 1570
rect 2032 1622 2182 1624
rect 2032 1570 2038 1622
rect 2090 1570 2124 1622
rect 2176 1570 2182 1622
rect 2032 1568 2182 1570
rect 2548 1622 2700 1624
rect 2548 1570 2554 1622
rect 2606 1613 2700 1622
rect 2606 1579 2649 1613
rect 2683 1579 2700 1613
rect 2606 1570 2700 1579
rect 2548 1568 2700 1570
rect 482 1538 806 1540
rect 482 1529 748 1538
rect 482 1495 499 1529
rect 533 1495 748 1529
rect 482 1486 748 1495
rect 800 1486 806 1538
rect 482 1484 806 1486
rect 2116 1538 2354 1540
rect 2116 1529 2296 1538
rect 2116 1495 2133 1529
rect 2167 1495 2296 1529
rect 2116 1486 2296 1495
rect 2348 1486 2354 1538
rect 2116 1484 2354 1486
rect 226 1454 290 1456
rect 226 1402 232 1454
rect 284 1402 290 1454
rect 226 1400 290 1402
rect 1978 1445 2184 1456
rect 1978 1411 2133 1445
rect 2167 1411 2184 1445
rect 1978 1400 2184 1411
rect 2548 1454 2698 1456
rect 2548 1402 2554 1454
rect 2606 1402 2640 1454
rect 2692 1402 2698 1454
rect 2548 1400 2698 1402
rect 828 1370 892 1372
rect 828 1318 834 1370
rect 886 1318 892 1370
rect 828 1316 892 1318
rect 946 1361 1238 1372
rect 946 1327 1187 1361
rect 1221 1327 1238 1361
rect 946 1316 1238 1327
rect 1170 1286 1494 1288
rect 1170 1277 1436 1286
rect 1170 1243 1187 1277
rect 1221 1243 1436 1277
rect 1170 1234 1436 1243
rect 1488 1234 1494 1286
rect 1170 1232 1494 1234
rect 416 512 454 602
rect 828 110 978 112
rect 828 58 834 110
rect 886 58 920 110
rect 972 58 978 110
rect 828 56 978 58
rect 1256 26 1324 28
rect 1256 -26 1264 26
rect 1316 -26 1324 26
rect 1256 -28 1324 -26
rect 2632 26 2700 28
rect 2632 -26 2640 26
rect 2692 -26 2700 26
rect 2632 -28 2700 -26
<< via1 >>
rect 318 2830 370 2882
rect 834 2830 886 2882
rect 1350 1738 1402 1790
rect 232 1654 284 1706
rect 834 1570 886 1622
rect 2038 1570 2090 1622
rect 2124 1570 2176 1622
rect 2554 1570 2606 1622
rect 748 1486 800 1538
rect 2296 1486 2348 1538
rect 232 1402 284 1454
rect 2554 1402 2606 1454
rect 2640 1402 2692 1454
rect 834 1318 886 1370
rect 1436 1234 1488 1286
rect 834 58 886 110
rect 920 58 972 110
rect 1264 17 1316 26
rect 1264 -17 1273 17
rect 1273 -17 1307 17
rect 1307 -17 1316 17
rect 1264 -26 1316 -17
rect 2640 17 2692 26
rect 2640 -17 2649 17
rect 2649 -17 2683 17
rect 2683 -17 2692 17
rect 2640 -26 2692 -17
<< metal2 >>
rect 316 2882 372 2888
rect 316 2830 318 2882
rect 370 2830 372 2882
rect 144 1792 200 1801
rect 144 1344 200 1736
rect 316 1792 372 2830
rect 316 1727 372 1736
rect 832 2882 888 2888
rect 832 2830 834 2882
rect 886 2830 888 2882
rect 832 1792 888 2830
rect 832 1727 888 1736
rect 1262 1792 1318 1801
rect 230 1706 286 1712
rect 230 1654 232 1706
rect 284 1654 286 1706
rect 230 1454 286 1654
rect 832 1622 888 1628
rect 832 1570 834 1622
rect 886 1570 888 1622
rect 230 1402 232 1454
rect 284 1402 286 1454
rect 746 1538 802 1544
rect 746 1486 748 1538
rect 800 1486 802 1538
rect 746 1428 802 1486
rect 230 1396 286 1402
rect 832 1370 888 1570
rect 832 1318 834 1370
rect 886 1318 888 1370
rect 832 1312 888 1318
rect 1262 1288 1318 1736
rect 1348 1790 1404 1796
rect 1348 1738 1350 1790
rect 1402 1738 1404 1790
rect 1348 1732 1404 1738
rect 2638 1792 2694 1801
rect 2036 1622 2092 1680
rect 2036 1570 2038 1622
rect 2090 1570 2092 1622
rect 2036 1564 2092 1570
rect 2122 1622 2178 1628
rect 2122 1570 2124 1622
rect 2176 1570 2178 1622
rect 1262 1223 1318 1232
rect 1348 1288 1404 1297
rect 1348 1223 1404 1232
rect 1434 1286 1490 1292
rect 1434 1234 1436 1286
rect 1488 1234 1490 1286
rect 1434 1228 1490 1234
rect 2036 1288 2092 1297
rect 2036 1223 2092 1232
rect 832 110 888 116
rect 832 58 834 110
rect 886 58 888 110
rect 832 28 888 58
rect 918 110 974 168
rect 918 58 920 110
rect 972 58 974 110
rect 918 52 974 58
rect 832 -37 888 -28
rect 1262 28 1318 48
rect 1262 -37 1318 -28
rect 2122 28 2178 1570
rect 2552 1622 2608 1680
rect 2552 1570 2554 1622
rect 2606 1570 2608 1622
rect 2552 1564 2608 1570
rect 2294 1538 2350 1544
rect 2294 1486 2296 1538
rect 2348 1486 2350 1538
rect 2294 1480 2350 1486
rect 2552 1454 2608 1460
rect 2552 1402 2554 1454
rect 2606 1402 2608 1454
rect 2552 1344 2608 1402
rect 2638 1454 2694 1736
rect 2638 1402 2640 1454
rect 2692 1402 2694 1454
rect 2638 1396 2694 1402
rect 2122 -37 2178 -28
rect 2638 28 2694 48
rect 2638 -37 2694 -28
<< via2 >>
rect 144 1736 200 1792
rect 316 1736 372 1792
rect 832 1736 888 1792
rect 1262 1736 1318 1792
rect 2638 1736 2694 1792
rect 1262 1232 1318 1288
rect 1348 1232 1404 1288
rect 2036 1232 2092 1288
rect 832 -28 888 28
rect 1262 26 1318 28
rect 1262 -26 1264 26
rect 1264 -26 1316 26
rect 1316 -26 1318 26
rect 1262 -28 1318 -26
rect 2122 -28 2178 28
rect 2638 26 2694 28
rect 2638 -26 2640 26
rect 2640 -26 2692 26
rect 2692 -26 2694 26
rect 2638 -28 2694 -26
<< metal3 >>
rect -80 1796 2832 1844
rect -80 1792 2040 1796
rect -80 1736 144 1792
rect 200 1736 316 1792
rect 372 1736 832 1792
rect 888 1736 1262 1792
rect 1318 1736 2040 1792
rect -80 1732 2040 1736
rect 2104 1732 2336 1796
rect 2400 1792 2832 1796
rect 2400 1736 2638 1792
rect 2694 1736 2832 1792
rect 2400 1732 2832 1736
rect -80 1684 2832 1732
rect 1257 1288 1409 1340
rect 1257 1232 1262 1288
rect 1318 1232 1348 1288
rect 1404 1232 1409 1288
rect 1257 1180 1409 1232
rect 2031 1292 2105 1340
rect 2031 1288 2040 1292
rect 2031 1232 2036 1288
rect 2031 1228 2040 1232
rect 2104 1228 2105 1292
rect 2031 1180 2105 1228
rect -80 32 2832 80
rect -80 -32 -32 32
rect 32 28 2832 32
rect 32 -28 832 28
rect 888 -28 1262 28
rect 1318 -28 2122 28
rect 2178 -28 2638 28
rect 2694 -28 2832 28
rect 32 -32 2832 -28
rect -80 -80 2832 -32
<< via3 >>
rect 2040 1732 2104 1796
rect 2336 1732 2400 1796
rect 2040 1288 2104 1292
rect 2040 1232 2092 1288
rect 2092 1232 2104 1288
rect 2040 1228 2104 1232
rect -32 -32 32 32
<< metal4 >>
rect -118 32 118 1882
rect 1954 1796 2190 1797
rect 1954 1732 2040 1796
rect 2104 1732 2190 1796
rect 1954 1292 2190 1732
rect 1954 1228 2040 1292
rect 2104 1228 2190 1292
rect 1954 1227 2190 1228
rect 2250 1796 2486 1882
rect 2250 1732 2336 1796
rect 2400 1732 2486 1796
rect -118 -32 -32 32
rect 32 -32 118 32
rect -118 -118 118 -32
rect 2250 -118 2486 1732
use INV_72761973_PG0_0_0_1678373049  INV_72761973_PG0_0_0_1678373049_0
timestamp 1678373424
transform 1 0 2236 0 1 0
box 0 30 516 3024
use NMOS_4T_17534534_X1_Y1_1678373051  NMOS_4T_17534534_X1_Y1_1678373051_0
timestamp 1678373424
transform -1 0 1118 0 1 1512
box 52 56 395 1482
use NMOS_4T_17534534_X1_Y1_1678373051  NMOS_4T_17534534_X1_Y1_1678373051_1
timestamp 1678373424
transform -1 0 602 0 1 1512
box 52 56 395 1482
use NMOS_S_48172527_X1_Y1_1678373052  NMOS_S_48172527_X1_Y1_1678373052_0
timestamp 1678375764
transform -1 0 516 0 -1 1512
box 52 56 395 1482
use SCM_PMOS_98301772_X1_Y1_1678373053  SCM_PMOS_98301772_X1_Y1_1678373053_0
timestamp 1678373424
transform 1 0 516 0 -1 1512
box 0 0 688 1512
use STAGE2_INV_89790208_PG0_0_0_1678373050  STAGE2_INV_89790208_PG0_0_0_1678373050_0
timestamp 1678373424
transform -1 0 2236 0 1 0
box 0 30 1032 3024
<< labels >>
flabel metal1 s 2408 1428 2408 1428 0 FreeSerif 0 0 0 0 OUT
port 1 nsew
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
port 3 nsew
rlabel metal1 434 532 434 532 1 BIAS
port 6 n
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
port 2 nsew
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
rlabel metal1 1036 2478 1036 2478 1 INP
port 4 n
<< end >>
