magic
tech sky130A
magscale 1 2
timestamp 1678376823
<< error_p >>
rect 1204 1680 1458 1766
rect 1036 1512 1458 1680
rect 2004 1568 2012 1624
rect 2032 1568 2040 1624
rect 2520 1568 2528 1624
rect 2548 1568 2556 1624
rect 2520 1400 2528 1456
rect 2548 1400 2556 1456
<< nwell >>
rect 1204 1512 2752 3024
rect 516 0 1204 1512
<< pwell >>
rect 301 2718 387 2994
rect 817 2718 903 2994
rect 207 1969 481 2189
rect 723 1969 997 2189
rect 121 835 395 1055
rect 215 30 301 306
rect 1325 835 1599 1055
rect 1841 835 2115 1055
rect 2357 835 2631 1055
rect 1419 30 1505 306
rect 1935 30 2021 306
rect 2451 30 2537 306
<< nmos >>
rect 286 1995 316 2163
rect 372 1995 402 2163
rect 802 1995 832 2163
rect 888 1995 918 2163
rect 200 861 230 1029
rect 286 861 316 1029
rect 1404 861 1434 1029
rect 1490 861 1520 1029
rect 1920 861 1950 1029
rect 2006 861 2036 1029
rect 2436 861 2466 1029
rect 2522 861 2552 1029
<< pmos >>
rect 1404 1995 1434 2163
rect 1490 1995 1520 2163
rect 1920 1995 1950 2163
rect 2006 1995 2036 2163
rect 2436 1995 2466 2163
rect 2522 1995 2552 2163
rect 716 861 746 1029
rect 802 861 832 1029
rect 888 861 918 1029
rect 974 861 1004 1029
<< ndiff >>
rect 233 2113 286 2163
rect 233 2079 241 2113
rect 275 2079 286 2113
rect 233 2045 286 2079
rect 233 2011 241 2045
rect 275 2011 286 2045
rect 233 1995 286 2011
rect 316 2113 372 2163
rect 316 2079 327 2113
rect 361 2079 372 2113
rect 316 2045 372 2079
rect 316 2011 327 2045
rect 361 2011 372 2045
rect 316 1995 372 2011
rect 402 2113 455 2163
rect 402 2079 413 2113
rect 447 2079 455 2113
rect 402 2045 455 2079
rect 402 2011 413 2045
rect 447 2011 455 2045
rect 402 1995 455 2011
rect 749 2113 802 2163
rect 749 2079 757 2113
rect 791 2079 802 2113
rect 749 2045 802 2079
rect 749 2011 757 2045
rect 791 2011 802 2045
rect 749 1995 802 2011
rect 832 2113 888 2163
rect 832 2079 843 2113
rect 877 2079 888 2113
rect 832 2045 888 2079
rect 832 2011 843 2045
rect 877 2011 888 2045
rect 832 1995 888 2011
rect 918 2113 971 2163
rect 918 2079 929 2113
rect 963 2079 971 2113
rect 918 2045 971 2079
rect 918 2011 929 2045
rect 963 2011 971 2045
rect 918 1995 971 2011
rect 147 1013 200 1029
rect 147 979 155 1013
rect 189 979 200 1013
rect 147 945 200 979
rect 147 911 155 945
rect 189 911 200 945
rect 147 861 200 911
rect 230 1013 286 1029
rect 230 979 241 1013
rect 275 979 286 1013
rect 230 945 286 979
rect 230 911 241 945
rect 275 911 286 945
rect 230 861 286 911
rect 316 1013 369 1029
rect 316 979 327 1013
rect 361 979 369 1013
rect 316 945 369 979
rect 316 911 327 945
rect 361 911 369 945
rect 316 861 369 911
rect 1351 1013 1404 1029
rect 1351 979 1359 1013
rect 1393 979 1404 1013
rect 1351 945 1404 979
rect 1351 911 1359 945
rect 1393 911 1404 945
rect 1351 861 1404 911
rect 1434 1013 1490 1029
rect 1434 979 1445 1013
rect 1479 979 1490 1013
rect 1434 945 1490 979
rect 1434 911 1445 945
rect 1479 911 1490 945
rect 1434 861 1490 911
rect 1520 1013 1573 1029
rect 1520 979 1531 1013
rect 1565 979 1573 1013
rect 1520 945 1573 979
rect 1520 911 1531 945
rect 1565 911 1573 945
rect 1520 861 1573 911
rect 1867 1013 1920 1029
rect 1867 979 1875 1013
rect 1909 979 1920 1013
rect 1867 945 1920 979
rect 1867 911 1875 945
rect 1909 911 1920 945
rect 1867 861 1920 911
rect 1950 1013 2006 1029
rect 1950 979 1961 1013
rect 1995 979 2006 1013
rect 1950 945 2006 979
rect 1950 911 1961 945
rect 1995 911 2006 945
rect 1950 861 2006 911
rect 2036 1013 2089 1029
rect 2036 979 2047 1013
rect 2081 979 2089 1013
rect 2036 945 2089 979
rect 2036 911 2047 945
rect 2081 911 2089 945
rect 2036 861 2089 911
rect 2383 1013 2436 1029
rect 2383 979 2391 1013
rect 2425 979 2436 1013
rect 2383 945 2436 979
rect 2383 911 2391 945
rect 2425 911 2436 945
rect 2383 861 2436 911
rect 2466 1013 2522 1029
rect 2466 979 2477 1013
rect 2511 979 2522 1013
rect 2466 945 2522 979
rect 2466 911 2477 945
rect 2511 911 2522 945
rect 2466 861 2522 911
rect 2552 1013 2605 1029
rect 2552 979 2563 1013
rect 2597 979 2605 1013
rect 2552 945 2605 979
rect 2552 911 2563 945
rect 2597 911 2605 945
rect 2552 861 2605 911
<< pdiff >>
rect 1351 2113 1404 2163
rect 1351 2079 1359 2113
rect 1393 2079 1404 2113
rect 1351 2045 1404 2079
rect 1351 2011 1359 2045
rect 1393 2011 1404 2045
rect 1351 1995 1404 2011
rect 1434 2113 1490 2163
rect 1434 2079 1445 2113
rect 1479 2079 1490 2113
rect 1434 2045 1490 2079
rect 1434 2011 1445 2045
rect 1479 2011 1490 2045
rect 1434 1995 1490 2011
rect 1520 2113 1573 2163
rect 1520 2079 1531 2113
rect 1565 2079 1573 2113
rect 1520 2045 1573 2079
rect 1520 2011 1531 2045
rect 1565 2011 1573 2045
rect 1520 1995 1573 2011
rect 1867 2113 1920 2163
rect 1867 2079 1875 2113
rect 1909 2079 1920 2113
rect 1867 2045 1920 2079
rect 1867 2011 1875 2045
rect 1909 2011 1920 2045
rect 1867 1995 1920 2011
rect 1950 2113 2006 2163
rect 1950 2079 1961 2113
rect 1995 2079 2006 2113
rect 1950 2045 2006 2079
rect 1950 2011 1961 2045
rect 1995 2011 2006 2045
rect 1950 1995 2006 2011
rect 2036 2113 2089 2163
rect 2036 2079 2047 2113
rect 2081 2079 2089 2113
rect 2036 2045 2089 2079
rect 2036 2011 2047 2045
rect 2081 2011 2089 2045
rect 2036 1995 2089 2011
rect 2383 2113 2436 2163
rect 2383 2079 2391 2113
rect 2425 2079 2436 2113
rect 2383 2045 2436 2079
rect 2383 2011 2391 2045
rect 2425 2011 2436 2045
rect 2383 1995 2436 2011
rect 2466 2113 2522 2163
rect 2466 2079 2477 2113
rect 2511 2079 2522 2113
rect 2466 2045 2522 2079
rect 2466 2011 2477 2045
rect 2511 2011 2522 2045
rect 2466 1995 2522 2011
rect 2552 2113 2605 2163
rect 2552 2079 2563 2113
rect 2597 2079 2605 2113
rect 2552 2045 2605 2079
rect 2552 2011 2563 2045
rect 2597 2011 2605 2045
rect 2552 1995 2605 2011
rect 663 1013 716 1029
rect 663 979 671 1013
rect 705 979 716 1013
rect 663 945 716 979
rect 663 911 671 945
rect 705 911 716 945
rect 663 861 716 911
rect 746 1013 802 1029
rect 746 979 757 1013
rect 791 979 802 1013
rect 746 945 802 979
rect 746 911 757 945
rect 791 911 802 945
rect 746 861 802 911
rect 832 1013 888 1029
rect 832 979 843 1013
rect 877 979 888 1013
rect 832 945 888 979
rect 832 911 843 945
rect 877 911 888 945
rect 832 861 888 911
rect 918 1013 974 1029
rect 918 979 929 1013
rect 963 979 974 1013
rect 918 945 974 979
rect 918 911 929 945
rect 963 911 974 945
rect 918 861 974 911
rect 1004 1013 1057 1029
rect 1004 979 1015 1013
rect 1049 979 1057 1013
rect 1004 945 1057 979
rect 1004 911 1015 945
rect 1049 911 1057 945
rect 1004 861 1057 911
<< ndiffc >>
rect 241 2079 275 2113
rect 241 2011 275 2045
rect 327 2079 361 2113
rect 327 2011 361 2045
rect 413 2079 447 2113
rect 413 2011 447 2045
rect 757 2079 791 2113
rect 757 2011 791 2045
rect 843 2079 877 2113
rect 843 2011 877 2045
rect 929 2079 963 2113
rect 929 2011 963 2045
rect 155 979 189 1013
rect 155 911 189 945
rect 241 979 275 1013
rect 241 911 275 945
rect 327 979 361 1013
rect 327 911 361 945
rect 1359 979 1393 1013
rect 1359 911 1393 945
rect 1445 979 1479 1013
rect 1445 911 1479 945
rect 1531 979 1565 1013
rect 1531 911 1565 945
rect 1875 979 1909 1013
rect 1875 911 1909 945
rect 1961 979 1995 1013
rect 1961 911 1995 945
rect 2047 979 2081 1013
rect 2047 911 2081 945
rect 2391 979 2425 1013
rect 2391 911 2425 945
rect 2477 979 2511 1013
rect 2477 911 2511 945
rect 2563 979 2597 1013
rect 2563 911 2597 945
<< pdiffc >>
rect 1359 2079 1393 2113
rect 1359 2011 1393 2045
rect 1445 2079 1479 2113
rect 1445 2011 1479 2045
rect 1531 2079 1565 2113
rect 1531 2011 1565 2045
rect 1875 2079 1909 2113
rect 1875 2011 1909 2045
rect 1961 2079 1995 2113
rect 1961 2011 1995 2045
rect 2047 2079 2081 2113
rect 2047 2011 2081 2045
rect 2391 2079 2425 2113
rect 2391 2011 2425 2045
rect 2477 2079 2511 2113
rect 2477 2011 2511 2045
rect 2563 2079 2597 2113
rect 2563 2011 2597 2045
rect 671 979 705 1013
rect 671 911 705 945
rect 757 979 791 1013
rect 757 911 791 945
rect 843 979 877 1013
rect 843 911 877 945
rect 929 979 963 1013
rect 929 911 963 945
rect 1015 979 1049 1013
rect 1015 911 1049 945
<< psubdiff >>
rect 327 2873 361 2968
rect 327 2744 361 2839
rect 843 2873 877 2968
rect 843 2744 877 2839
rect 241 185 275 280
rect 241 56 275 151
rect 1445 185 1479 280
rect 1445 56 1479 151
rect 1961 185 1995 280
rect 1961 56 1995 151
rect 2477 185 2511 280
rect 2477 56 2511 151
<< nsubdiff >>
rect 1445 2873 1479 2968
rect 1445 2744 1479 2839
rect 1961 2873 1995 2968
rect 1961 2744 1995 2839
rect 2477 2873 2511 2968
rect 2477 2744 2511 2839
rect 757 185 791 280
rect 757 56 791 151
rect 929 185 963 280
rect 929 56 963 151
<< psubdiffcont >>
rect 327 2839 361 2873
rect 843 2839 877 2873
rect 241 151 275 185
rect 1445 151 1479 185
rect 1961 151 1995 185
rect 2477 151 2511 185
<< nsubdiffcont >>
rect 1445 2839 1479 2873
rect 1961 2839 1995 2873
rect 2477 2839 2511 2873
rect 757 151 791 185
rect 929 151 963 185
<< poly >>
rect 286 2453 402 2463
rect 286 2419 327 2453
rect 361 2419 402 2453
rect 286 2409 402 2419
rect 286 2163 316 2409
rect 372 2163 402 2409
rect 802 2453 918 2463
rect 802 2419 843 2453
rect 877 2419 918 2453
rect 802 2409 918 2419
rect 802 2163 832 2409
rect 888 2163 918 2409
rect 1404 2453 1520 2463
rect 1404 2419 1445 2453
rect 1479 2419 1520 2453
rect 1404 2409 1520 2419
rect 1404 2163 1434 2409
rect 1490 2163 1520 2409
rect 1920 2453 2036 2463
rect 1920 2419 1961 2453
rect 1995 2419 2036 2453
rect 1920 2409 2036 2419
rect 1920 2163 1950 2409
rect 2006 2163 2036 2409
rect 2436 2453 2552 2463
rect 2436 2419 2477 2453
rect 2511 2419 2552 2453
rect 2436 2409 2552 2419
rect 2436 2163 2466 2409
rect 2522 2163 2552 2409
rect 286 1764 316 1995
rect 372 1764 402 1995
rect 802 1764 832 1995
rect 888 1764 918 1995
rect 1404 1764 1434 1995
rect 1490 1764 1520 1995
rect 1920 1764 1950 1995
rect 2006 1764 2036 1995
rect 2436 1764 2466 1995
rect 2522 1764 2552 1995
rect 200 1029 230 1260
rect 286 1029 316 1260
rect 716 1029 746 1260
rect 802 1029 832 1260
rect 888 1029 918 1260
rect 974 1029 1004 1260
rect 1404 1029 1434 1260
rect 1490 1029 1520 1260
rect 1920 1029 1950 1260
rect 2006 1029 2036 1260
rect 2436 1029 2466 1260
rect 2522 1029 2552 1260
rect 200 615 230 861
rect 286 615 316 861
rect 200 605 316 615
rect 200 571 241 605
rect 275 571 316 605
rect 200 561 316 571
rect 716 615 746 861
rect 802 615 832 861
rect 716 605 832 615
rect 716 571 757 605
rect 791 571 832 605
rect 716 561 832 571
rect 888 615 918 861
rect 974 615 1004 861
rect 888 605 1004 615
rect 888 571 929 605
rect 963 571 1004 605
rect 888 561 1004 571
rect 1404 615 1434 861
rect 1490 615 1520 861
rect 1404 605 1520 615
rect 1404 571 1445 605
rect 1479 571 1520 605
rect 1404 561 1520 571
rect 1920 615 1950 861
rect 2006 615 2036 861
rect 1920 605 2036 615
rect 1920 571 1961 605
rect 1995 571 2036 605
rect 1920 561 2036 571
rect 2436 615 2466 861
rect 2522 615 2552 861
rect 2436 605 2552 615
rect 2436 571 2477 605
rect 2511 571 2552 605
rect 2436 561 2552 571
<< polycont >>
rect 327 2419 361 2453
rect 843 2419 877 2453
rect 1445 2419 1479 2453
rect 1961 2419 1995 2453
rect 2477 2419 2511 2453
rect 241 571 275 605
rect 757 571 791 605
rect 929 571 963 605
rect 1445 571 1479 605
rect 1961 571 1995 605
rect 2477 571 2511 605
<< locali >>
rect 319 2873 369 2957
rect 319 2839 327 2873
rect 361 2839 369 2873
rect 319 2755 369 2839
rect 835 2873 885 2957
rect 835 2839 843 2873
rect 877 2839 885 2873
rect 835 2755 885 2839
rect 1437 2873 1487 2957
rect 1437 2839 1445 2873
rect 1479 2839 1487 2873
rect 1437 2755 1487 2839
rect 1953 2873 2003 2957
rect 1953 2839 1961 2873
rect 1995 2839 2003 2873
rect 1953 2755 2003 2839
rect 2469 2873 2519 2957
rect 2469 2839 2477 2873
rect 2511 2839 2519 2873
rect 2469 2755 2519 2839
rect 319 2453 369 2537
rect 319 2419 327 2453
rect 361 2419 369 2453
rect 319 2335 369 2419
rect 835 2453 885 2537
rect 835 2419 843 2453
rect 877 2419 885 2453
rect 835 2335 885 2419
rect 1437 2453 1487 2537
rect 1953 2453 2003 2537
rect 1437 2419 1445 2453
rect 1479 2419 1487 2453
rect 1437 2335 1487 2419
rect 1781 2419 1789 2453
rect 1823 2419 1831 2453
rect 1781 2369 1831 2419
rect 1609 2335 1617 2369
rect 1651 2335 1659 2369
rect 1781 2335 1789 2369
rect 1823 2335 1831 2369
rect 1953 2419 1961 2453
rect 1995 2419 2003 2453
rect 1953 2335 2003 2419
rect 2469 2453 2519 2537
rect 2469 2419 2477 2453
rect 2511 2419 2519 2453
rect 2469 2335 2519 2419
rect 233 2113 283 2285
rect 233 2079 241 2113
rect 275 2079 283 2113
rect 233 2045 283 2079
rect 233 2011 241 2045
rect 275 2011 283 2045
rect 233 1697 283 2011
rect 233 1663 241 1697
rect 275 1663 283 1697
rect 233 1579 283 1663
rect 319 2113 369 2285
rect 319 2079 327 2113
rect 361 2079 369 2113
rect 319 2045 369 2079
rect 319 2011 327 2045
rect 361 2011 369 2045
rect 319 1613 369 2011
rect 319 1579 327 1613
rect 361 1579 369 1613
rect 405 2113 455 2285
rect 405 2079 413 2113
rect 447 2079 455 2113
rect 405 2045 455 2079
rect 405 2011 413 2045
rect 447 2011 455 2045
rect 405 1697 455 2011
rect 405 1663 413 1697
rect 447 1663 455 1697
rect 405 1579 455 1663
rect 749 2113 799 2285
rect 749 2079 757 2113
rect 791 2079 799 2113
rect 749 2045 799 2079
rect 749 2011 757 2045
rect 791 2011 799 2045
rect 749 1697 799 2011
rect 749 1663 757 1697
rect 791 1663 799 1697
rect 491 1579 499 1613
rect 533 1579 541 1613
rect 749 1579 799 1663
rect 835 2113 885 2285
rect 835 2079 843 2113
rect 877 2079 885 2113
rect 835 2045 885 2079
rect 835 2011 843 2045
rect 877 2011 885 2045
rect 835 1613 885 2011
rect 835 1579 843 1613
rect 877 1579 885 1613
rect 921 2113 971 2285
rect 921 2079 929 2113
rect 963 2079 971 2113
rect 921 2045 971 2079
rect 921 2011 929 2045
rect 963 2011 971 2045
rect 921 1697 971 2011
rect 1351 2113 1401 2285
rect 1351 2079 1359 2113
rect 1393 2079 1401 2113
rect 1351 2045 1401 2079
rect 1351 2011 1359 2045
rect 1393 2011 1401 2045
rect 921 1663 929 1697
rect 963 1663 971 1697
rect 921 1579 971 1663
rect 1265 1747 1273 1781
rect 1307 1747 1315 1781
rect 491 1529 541 1579
rect 491 1495 499 1529
rect 533 1495 541 1529
rect 147 1361 197 1445
rect 147 1327 155 1361
rect 189 1327 197 1361
rect 147 1013 197 1327
rect 147 979 155 1013
rect 189 979 197 1013
rect 147 945 197 979
rect 147 911 155 945
rect 189 911 197 945
rect 147 739 197 911
rect 233 1411 241 1445
rect 275 1411 283 1445
rect 233 1013 283 1411
rect 233 979 241 1013
rect 275 979 283 1013
rect 233 945 283 979
rect 233 911 241 945
rect 275 911 283 945
rect 233 739 283 911
rect 319 1361 369 1445
rect 319 1327 327 1361
rect 361 1327 369 1361
rect 319 1013 369 1327
rect 319 979 327 1013
rect 361 979 369 1013
rect 319 945 369 979
rect 319 911 327 945
rect 361 911 369 945
rect 319 739 369 911
rect 663 1277 713 1445
rect 663 1243 671 1277
rect 705 1243 713 1277
rect 663 1013 713 1243
rect 663 979 671 1013
rect 705 979 713 1013
rect 663 945 713 979
rect 663 911 671 945
rect 705 911 713 945
rect 663 739 713 911
rect 749 1411 757 1445
rect 791 1411 799 1445
rect 749 1013 799 1411
rect 749 979 757 1013
rect 791 979 799 1013
rect 749 945 799 979
rect 749 911 757 945
rect 791 911 799 945
rect 749 739 799 911
rect 835 1277 885 1445
rect 835 1243 843 1277
rect 877 1243 885 1277
rect 835 1013 885 1243
rect 835 979 843 1013
rect 877 979 885 1013
rect 835 945 885 979
rect 835 911 843 945
rect 877 911 885 945
rect 835 739 885 911
rect 921 1361 971 1445
rect 921 1327 929 1361
rect 963 1327 971 1361
rect 921 1013 971 1327
rect 921 979 929 1013
rect 963 979 971 1013
rect 921 945 971 979
rect 921 911 929 945
rect 963 911 971 945
rect 921 739 971 911
rect 1007 1277 1057 1445
rect 1007 1243 1015 1277
rect 1049 1243 1057 1277
rect 1179 1327 1187 1361
rect 1221 1327 1229 1361
rect 1179 1277 1229 1327
rect 1179 1243 1187 1277
rect 1221 1243 1229 1277
rect 1007 1013 1057 1243
rect 1007 979 1015 1013
rect 1049 979 1057 1013
rect 1007 945 1057 979
rect 1007 911 1015 945
rect 1049 911 1057 945
rect 1007 739 1057 911
rect 233 605 283 689
rect 233 571 241 605
rect 275 571 283 605
rect 233 487 283 571
rect 749 605 799 689
rect 749 571 757 605
rect 791 571 799 605
rect 749 487 799 571
rect 921 605 971 689
rect 921 571 929 605
rect 963 571 971 605
rect 921 487 971 571
rect 233 185 283 269
rect 233 151 241 185
rect 275 151 283 185
rect 233 67 283 151
rect 749 185 799 269
rect 749 151 757 185
rect 791 151 799 185
rect 749 67 799 151
rect 921 185 971 269
rect 921 151 929 185
rect 963 151 971 185
rect 921 67 971 151
rect 1265 17 1315 1747
rect 1351 1697 1401 2011
rect 1351 1663 1359 1697
rect 1393 1663 1401 1697
rect 1351 1579 1401 1663
rect 1437 2113 1487 2285
rect 1437 2079 1445 2113
rect 1479 2079 1487 2113
rect 1437 2045 1487 2079
rect 1437 2011 1445 2045
rect 1479 2011 1487 2045
rect 1437 1613 1487 2011
rect 1437 1579 1445 1613
rect 1479 1579 1487 1613
rect 1523 2113 1573 2285
rect 1523 2079 1531 2113
rect 1565 2079 1573 2113
rect 1523 2045 1573 2079
rect 1523 2011 1531 2045
rect 1565 2011 1573 2045
rect 1523 1697 1573 2011
rect 1523 1663 1531 1697
rect 1565 1663 1573 1697
rect 1523 1579 1573 1663
rect 1609 1613 1659 2335
rect 1867 2113 1917 2285
rect 1867 2079 1875 2113
rect 1909 2079 1917 2113
rect 1867 2045 1917 2079
rect 1867 2011 1875 2045
rect 1909 2011 1917 2045
rect 1867 1697 1917 2011
rect 1867 1663 1875 1697
rect 1909 1663 1917 1697
rect 1609 1579 1617 1613
rect 1651 1579 1659 1613
rect 1609 1445 1659 1579
rect 1351 1361 1401 1445
rect 1351 1327 1359 1361
rect 1393 1327 1401 1361
rect 1351 1013 1401 1327
rect 1351 979 1359 1013
rect 1393 979 1401 1013
rect 1351 945 1401 979
rect 1351 911 1359 945
rect 1393 911 1401 945
rect 1351 739 1401 911
rect 1437 1411 1445 1445
rect 1479 1411 1487 1445
rect 1437 1013 1487 1411
rect 1437 979 1445 1013
rect 1479 979 1487 1013
rect 1437 945 1487 979
rect 1437 911 1445 945
rect 1479 911 1487 945
rect 1437 739 1487 911
rect 1523 1361 1573 1445
rect 1523 1327 1531 1361
rect 1565 1327 1573 1361
rect 1523 1013 1573 1327
rect 1609 1411 1617 1445
rect 1651 1411 1659 1445
rect 1781 1579 1789 1613
rect 1823 1579 1831 1613
rect 1867 1579 1917 1663
rect 1953 2113 2003 2285
rect 1953 2079 1961 2113
rect 1995 2079 2003 2113
rect 1953 2045 2003 2079
rect 1953 2011 1961 2045
rect 1995 2011 2003 2045
rect 1953 1613 2003 2011
rect 1953 1579 1961 1613
rect 1995 1579 2003 1613
rect 2039 2113 2089 2285
rect 2039 2079 2047 2113
rect 2081 2079 2089 2113
rect 2039 2045 2089 2079
rect 2039 2011 2047 2045
rect 2081 2011 2089 2045
rect 2039 1697 2089 2011
rect 2039 1663 2047 1697
rect 2081 1663 2089 1697
rect 2039 1579 2089 1663
rect 2383 2113 2433 2285
rect 2383 2079 2391 2113
rect 2425 2079 2433 2113
rect 2383 2045 2433 2079
rect 2383 2011 2391 2045
rect 2425 2011 2433 2045
rect 2383 1697 2433 2011
rect 2383 1663 2391 1697
rect 2425 1663 2433 1697
rect 2297 1579 2305 1613
rect 2339 1579 2347 1613
rect 2383 1579 2433 1663
rect 2469 2113 2519 2285
rect 2469 2079 2477 2113
rect 2511 2079 2519 2113
rect 2469 2045 2519 2079
rect 2469 2011 2477 2045
rect 2511 2011 2519 2045
rect 2469 1613 2519 2011
rect 2469 1579 2477 1613
rect 2511 1579 2519 1613
rect 2555 2113 2605 2285
rect 2555 2079 2563 2113
rect 2597 2079 2605 2113
rect 2555 2045 2605 2079
rect 2555 2011 2563 2045
rect 2597 2011 2605 2045
rect 2555 1697 2605 2011
rect 2555 1663 2563 1697
rect 2597 1663 2605 1697
rect 2555 1579 2605 1663
rect 2641 1579 2649 1613
rect 2683 1579 2691 1613
rect 1781 1445 1831 1579
rect 2125 1495 2133 1529
rect 2167 1495 2175 1529
rect 2125 1445 2175 1495
rect 1781 1411 1789 1445
rect 1823 1411 1831 1445
rect 1609 1277 1659 1411
rect 1867 1361 1917 1445
rect 1867 1327 1875 1361
rect 1909 1327 1917 1361
rect 1609 1243 1617 1277
rect 1651 1243 1659 1277
rect 1781 1243 1789 1277
rect 1823 1243 1831 1277
rect 1523 979 1531 1013
rect 1565 979 1573 1013
rect 1523 945 1573 979
rect 1523 911 1531 945
rect 1565 911 1573 945
rect 1523 739 1573 911
rect 1437 605 1487 689
rect 1437 571 1445 605
rect 1479 571 1487 605
rect 1781 605 1831 1243
rect 1867 1013 1917 1327
rect 1867 979 1875 1013
rect 1909 979 1917 1013
rect 1867 945 1917 979
rect 1867 911 1875 945
rect 1909 911 1917 945
rect 1867 739 1917 911
rect 1953 1411 1961 1445
rect 1995 1411 2003 1445
rect 1953 1013 2003 1411
rect 1953 979 1961 1013
rect 1995 979 2003 1013
rect 1953 945 2003 979
rect 1953 911 1961 945
rect 1995 911 2003 945
rect 1953 739 2003 911
rect 2039 1361 2089 1445
rect 2125 1411 2133 1445
rect 2167 1411 2175 1445
rect 2297 1445 2347 1579
rect 2297 1411 2305 1445
rect 2339 1411 2347 1445
rect 2039 1327 2047 1361
rect 2081 1327 2089 1361
rect 2039 1013 2089 1327
rect 2039 979 2047 1013
rect 2081 979 2089 1013
rect 2039 945 2089 979
rect 2039 911 2047 945
rect 2081 911 2089 945
rect 2039 739 2089 911
rect 2383 1361 2433 1445
rect 2383 1327 2391 1361
rect 2425 1327 2433 1361
rect 2383 1013 2433 1327
rect 2383 979 2391 1013
rect 2425 979 2433 1013
rect 2383 945 2433 979
rect 2383 911 2391 945
rect 2425 911 2433 945
rect 2383 739 2433 911
rect 2469 1411 2477 1445
rect 2511 1411 2519 1445
rect 2469 1013 2519 1411
rect 2469 979 2477 1013
rect 2511 979 2519 1013
rect 2469 945 2519 979
rect 2469 911 2477 945
rect 2511 911 2519 945
rect 2469 739 2519 911
rect 2555 1361 2605 1445
rect 2555 1327 2563 1361
rect 2597 1327 2605 1361
rect 2555 1013 2605 1327
rect 2555 979 2563 1013
rect 2597 979 2605 1013
rect 2555 945 2605 979
rect 2555 911 2563 945
rect 2597 911 2605 945
rect 2555 739 2605 911
rect 1781 571 1789 605
rect 1823 571 1831 605
rect 1953 605 2003 689
rect 1953 571 1961 605
rect 1995 571 2003 605
rect 1437 487 1487 571
rect 1953 487 2003 571
rect 2469 605 2519 689
rect 2469 571 2477 605
rect 2511 571 2519 605
rect 2469 487 2519 571
rect 1437 185 1487 269
rect 1437 151 1445 185
rect 1479 151 1487 185
rect 1437 67 1487 151
rect 1953 185 2003 269
rect 1953 151 1961 185
rect 1995 151 2003 185
rect 1953 67 2003 151
rect 2469 185 2519 269
rect 2469 151 2477 185
rect 2511 151 2519 185
rect 2469 67 2519 151
rect 1265 -17 1273 17
rect 1307 -17 1315 17
rect 2641 17 2691 1579
rect 2641 -17 2649 17
rect 2683 -17 2691 17
<< viali >>
rect 327 2839 361 2873
rect 843 2839 877 2873
rect 1445 2839 1479 2873
rect 1961 2839 1995 2873
rect 2477 2839 2511 2873
rect 327 2419 361 2453
rect 843 2419 877 2453
rect 1445 2419 1479 2453
rect 1789 2419 1823 2453
rect 1617 2335 1651 2369
rect 1789 2335 1823 2369
rect 1961 2419 1995 2453
rect 2477 2419 2511 2453
rect 241 1663 275 1697
rect 327 1579 361 1613
rect 413 1663 447 1697
rect 757 1663 791 1697
rect 499 1579 533 1613
rect 843 1579 877 1613
rect 929 1663 963 1697
rect 1273 1747 1307 1781
rect 499 1495 533 1529
rect 155 1327 189 1361
rect 241 1411 275 1445
rect 327 1327 361 1361
rect 671 1243 705 1277
rect 757 1411 791 1445
rect 843 1243 877 1277
rect 929 1327 963 1361
rect 1015 1243 1049 1277
rect 1187 1327 1221 1361
rect 1187 1243 1221 1277
rect 241 571 275 605
rect 757 571 791 605
rect 929 571 963 605
rect 241 151 275 185
rect 757 151 791 185
rect 929 151 963 185
rect 1359 1663 1393 1697
rect 1445 1579 1479 1613
rect 1531 1663 1565 1697
rect 1875 1663 1909 1697
rect 1617 1579 1651 1613
rect 1359 1327 1393 1361
rect 1445 1411 1479 1445
rect 1531 1327 1565 1361
rect 1617 1411 1651 1445
rect 1789 1579 1823 1613
rect 1961 1579 1995 1613
rect 2047 1663 2081 1697
rect 2391 1663 2425 1697
rect 2305 1579 2339 1613
rect 2477 1579 2511 1613
rect 2563 1663 2597 1697
rect 2649 1579 2683 1613
rect 2133 1495 2167 1529
rect 1789 1411 1823 1445
rect 1875 1327 1909 1361
rect 1617 1243 1651 1277
rect 1789 1243 1823 1277
rect 1445 571 1479 605
rect 1961 1411 1995 1445
rect 2133 1411 2167 1445
rect 2305 1411 2339 1445
rect 2047 1327 2081 1361
rect 2391 1327 2425 1361
rect 2477 1411 2511 1445
rect 2563 1327 2597 1361
rect 1789 571 1823 605
rect 1961 571 1995 605
rect 2477 571 2511 605
rect 1445 151 1479 185
rect 1961 151 1995 185
rect 2477 151 2511 185
rect 1273 -17 1307 17
rect 2649 -17 2683 17
<< metal1 >>
rect 310 2882 550 2884
rect 310 2830 318 2882
rect 370 2830 550 2882
rect 310 2828 550 2830
rect 826 2882 1066 2884
rect 826 2830 834 2882
rect 886 2830 1066 2882
rect 826 2828 1066 2830
rect 1342 2882 1582 2884
rect 1342 2830 1350 2882
rect 1402 2873 1582 2882
rect 1402 2839 1445 2873
rect 1479 2839 1582 2873
rect 1402 2830 1582 2839
rect 1342 2828 1582 2830
rect 1858 2882 2098 2884
rect 1858 2873 2038 2882
rect 1858 2839 1961 2873
rect 1995 2839 2038 2873
rect 1858 2830 2038 2839
rect 2090 2830 2098 2882
rect 1858 2828 2098 2830
rect 2374 2882 2614 2884
rect 2374 2873 2554 2882
rect 2374 2839 2477 2873
rect 2511 2839 2554 2873
rect 2374 2830 2554 2839
rect 2606 2830 2614 2882
rect 2374 2828 2614 2830
rect 310 2453 550 2464
rect 310 2419 327 2453
rect 361 2419 550 2453
rect 310 2408 550 2419
rect 826 2453 1066 2464
rect 826 2419 843 2453
rect 877 2419 1066 2453
rect 826 2408 1066 2419
rect 1428 2462 1668 2464
rect 1428 2410 1436 2462
rect 1488 2410 1668 2462
rect 1428 2408 1668 2410
rect 1772 2453 2012 2464
rect 1772 2419 1789 2453
rect 1823 2419 1961 2453
rect 1995 2419 2012 2453
rect 1772 2408 2012 2419
rect 2288 2462 2528 2464
rect 2288 2410 2296 2462
rect 2348 2453 2528 2462
rect 2348 2419 2477 2453
rect 2511 2419 2528 2453
rect 2348 2410 2528 2419
rect 2288 2408 2528 2410
rect 1600 2369 1840 2380
rect 1600 2335 1617 2369
rect 1651 2335 1789 2369
rect 1823 2335 1840 2369
rect 1600 2324 1840 2335
rect 1256 1790 1408 1792
rect 1256 1781 1350 1790
rect 1256 1747 1273 1781
rect 1307 1747 1350 1781
rect 1256 1738 1350 1747
rect 1402 1738 1408 1790
rect 1256 1736 1408 1738
rect 224 1706 980 1708
rect 224 1654 232 1706
rect 284 1697 980 1706
rect 284 1663 413 1697
rect 447 1663 757 1697
rect 791 1663 929 1697
rect 963 1663 980 1697
rect 284 1654 980 1663
rect 224 1652 980 1654
rect 1342 1706 1582 1708
rect 1342 1654 1350 1706
rect 1402 1697 1582 1706
rect 1402 1663 1531 1697
rect 1565 1663 1582 1697
rect 1402 1654 1582 1663
rect 1342 1652 1582 1654
rect 1858 1706 2098 1708
rect 1858 1697 2038 1706
rect 1858 1663 1875 1697
rect 1909 1663 2038 1697
rect 1858 1654 2038 1663
rect 2090 1654 2098 1706
rect 1858 1652 2098 1654
rect 2374 1706 2614 1708
rect 2374 1697 2554 1706
rect 2374 1663 2391 1697
rect 2425 1663 2554 1697
rect 2374 1654 2554 1663
rect 2606 1654 2614 1706
rect 2374 1652 2614 1654
rect 310 1613 550 1624
rect 310 1579 327 1613
rect 361 1579 499 1613
rect 533 1579 550 1613
rect 310 1568 550 1579
rect 826 1622 1066 1624
rect 826 1570 834 1622
rect 886 1570 1066 1622
rect 826 1568 1066 1570
rect 1428 1613 1668 1624
rect 1428 1579 1445 1613
rect 1479 1579 1617 1613
rect 1651 1579 1668 1613
rect 1428 1568 1668 1579
rect 1772 1613 2012 1624
rect 1772 1579 1789 1613
rect 1823 1579 1961 1613
rect 1995 1579 2012 1613
rect 1772 1568 2012 1579
rect 2032 1622 2182 1624
rect 2032 1570 2038 1622
rect 2090 1570 2124 1622
rect 2176 1570 2182 1622
rect 2032 1568 2182 1570
rect 2288 1613 2528 1624
rect 2288 1579 2305 1613
rect 2339 1579 2477 1613
rect 2511 1579 2528 1613
rect 2288 1568 2528 1579
rect 2548 1622 2700 1624
rect 2548 1570 2554 1622
rect 2606 1613 2700 1622
rect 2606 1579 2649 1613
rect 2683 1579 2700 1613
rect 2606 1570 2700 1579
rect 2548 1568 2700 1570
rect 482 1538 806 1540
rect 482 1529 748 1538
rect 482 1495 499 1529
rect 533 1495 748 1529
rect 482 1486 748 1495
rect 800 1486 806 1538
rect 482 1484 806 1486
rect 2116 1538 2354 1540
rect 2116 1529 2296 1538
rect 2116 1495 2133 1529
rect 2167 1495 2296 1529
rect 2116 1486 2296 1495
rect 2348 1486 2354 1538
rect 2116 1484 2354 1486
rect 224 1454 464 1456
rect 224 1402 232 1454
rect 284 1402 464 1454
rect 224 1400 464 1402
rect 568 1454 808 1456
rect 568 1402 748 1454
rect 800 1402 808 1454
rect 568 1400 808 1402
rect 1428 1445 1668 1456
rect 1428 1411 1445 1445
rect 1479 1411 1617 1445
rect 1651 1411 1668 1445
rect 1428 1400 1668 1411
rect 1772 1445 2184 1456
rect 1772 1411 1789 1445
rect 1823 1411 1961 1445
rect 1995 1411 2133 1445
rect 2167 1411 2184 1445
rect 1772 1400 2184 1411
rect 2288 1445 2528 1456
rect 2288 1411 2305 1445
rect 2339 1411 2477 1445
rect 2511 1411 2528 1445
rect 2288 1400 2528 1411
rect 2548 1454 2698 1456
rect 2548 1402 2554 1454
rect 2606 1402 2640 1454
rect 2692 1402 2698 1454
rect 2548 1400 2698 1402
rect 138 1370 378 1372
rect 138 1318 146 1370
rect 198 1361 378 1370
rect 198 1327 327 1361
rect 361 1327 378 1361
rect 198 1318 378 1327
rect 138 1316 378 1318
rect 740 1370 1238 1372
rect 740 1318 834 1370
rect 886 1361 1238 1370
rect 886 1327 929 1361
rect 963 1327 1187 1361
rect 1221 1327 1238 1361
rect 886 1318 1238 1327
rect 740 1316 1238 1318
rect 1342 1370 1582 1372
rect 1342 1318 1350 1370
rect 1402 1361 1582 1370
rect 1402 1327 1531 1361
rect 1565 1327 1582 1361
rect 1402 1318 1582 1327
rect 1342 1316 1582 1318
rect 1858 1370 2098 1372
rect 1858 1361 2038 1370
rect 1858 1327 1875 1361
rect 1909 1327 2038 1361
rect 1858 1318 2038 1327
rect 2090 1318 2098 1370
rect 1858 1316 2098 1318
rect 2374 1370 2614 1372
rect 2374 1361 2554 1370
rect 2374 1327 2391 1361
rect 2425 1327 2554 1361
rect 2374 1318 2554 1327
rect 2606 1318 2614 1370
rect 2374 1316 2614 1318
rect 654 1286 1066 1288
rect 654 1277 920 1286
rect 654 1243 671 1277
rect 705 1243 843 1277
rect 877 1243 920 1277
rect 654 1234 920 1243
rect 972 1277 1066 1286
rect 972 1243 1015 1277
rect 1049 1243 1066 1277
rect 972 1234 1066 1243
rect 654 1232 1066 1234
rect 1170 1286 1494 1288
rect 1170 1277 1436 1286
rect 1170 1243 1187 1277
rect 1221 1243 1436 1277
rect 1170 1234 1436 1243
rect 1488 1234 1494 1286
rect 1170 1232 1494 1234
rect 1600 1277 1840 1288
rect 1600 1243 1617 1277
rect 1651 1243 1789 1277
rect 1823 1243 1840 1277
rect 1600 1232 1840 1243
rect 224 605 464 616
rect 224 571 241 605
rect 275 571 464 605
rect 224 560 464 571
rect 740 614 980 616
rect 740 562 748 614
rect 800 605 980 614
rect 800 571 929 605
rect 963 571 980 605
rect 800 562 980 571
rect 740 560 980 562
rect 1428 614 1668 616
rect 1428 562 1436 614
rect 1488 562 1668 614
rect 1428 560 1668 562
rect 1772 605 2012 616
rect 1772 571 1789 605
rect 1823 571 1961 605
rect 1995 571 2012 605
rect 1772 560 2012 571
rect 2288 614 2528 616
rect 2288 562 2296 614
rect 2348 605 2528 614
rect 2348 571 2477 605
rect 2511 571 2528 605
rect 2348 562 2528 571
rect 2288 560 2528 562
rect 138 194 378 196
rect 138 142 146 194
rect 198 185 378 194
rect 198 151 241 185
rect 275 151 378 185
rect 198 142 378 151
rect 138 140 378 142
rect 740 194 980 196
rect 740 185 920 194
rect 740 151 757 185
rect 791 151 920 185
rect 740 142 920 151
rect 972 142 980 194
rect 740 140 980 142
rect 1342 194 1582 196
rect 1342 142 1350 194
rect 1402 185 1582 194
rect 1402 151 1445 185
rect 1479 151 1582 185
rect 1402 142 1582 151
rect 1342 140 1582 142
rect 1858 194 2098 196
rect 1858 185 2038 194
rect 1858 151 1961 185
rect 1995 151 2038 185
rect 1858 142 2038 151
rect 2090 142 2098 194
rect 1858 140 2098 142
rect 2374 194 2614 196
rect 2374 185 2554 194
rect 2374 151 2477 185
rect 2511 151 2554 185
rect 2374 142 2554 151
rect 2606 142 2614 194
rect 2374 140 2614 142
rect 828 110 978 112
rect 828 58 834 110
rect 886 58 920 110
rect 972 58 978 110
rect 828 56 978 58
rect 1256 26 1324 28
rect 1256 -26 1264 26
rect 1316 -26 1324 26
rect 1256 -28 1324 -26
rect 2632 26 2700 28
rect 2632 -26 2640 26
rect 2692 -26 2700 26
rect 2632 -28 2700 -26
<< via1 >>
rect 318 2873 370 2882
rect 318 2839 327 2873
rect 327 2839 361 2873
rect 361 2839 370 2873
rect 318 2830 370 2839
rect 834 2873 886 2882
rect 834 2839 843 2873
rect 843 2839 877 2873
rect 877 2839 886 2873
rect 834 2830 886 2839
rect 1350 2830 1402 2882
rect 2038 2830 2090 2882
rect 2554 2830 2606 2882
rect 1436 2453 1488 2462
rect 1436 2419 1445 2453
rect 1445 2419 1479 2453
rect 1479 2419 1488 2453
rect 1436 2410 1488 2419
rect 2296 2410 2348 2462
rect 1350 1738 1402 1790
rect 232 1697 284 1706
rect 232 1663 241 1697
rect 241 1663 275 1697
rect 275 1663 284 1697
rect 232 1654 284 1663
rect 1350 1697 1402 1706
rect 1350 1663 1359 1697
rect 1359 1663 1393 1697
rect 1393 1663 1402 1697
rect 1350 1654 1402 1663
rect 2038 1697 2090 1706
rect 2038 1663 2047 1697
rect 2047 1663 2081 1697
rect 2081 1663 2090 1697
rect 2038 1654 2090 1663
rect 2554 1697 2606 1706
rect 2554 1663 2563 1697
rect 2563 1663 2597 1697
rect 2597 1663 2606 1697
rect 2554 1654 2606 1663
rect 834 1613 886 1622
rect 834 1579 843 1613
rect 843 1579 877 1613
rect 877 1579 886 1613
rect 834 1570 886 1579
rect 2038 1570 2090 1622
rect 2124 1570 2176 1622
rect 2554 1570 2606 1622
rect 748 1486 800 1538
rect 2296 1486 2348 1538
rect 232 1445 284 1454
rect 232 1411 241 1445
rect 241 1411 275 1445
rect 275 1411 284 1445
rect 232 1402 284 1411
rect 748 1445 800 1454
rect 748 1411 757 1445
rect 757 1411 791 1445
rect 791 1411 800 1445
rect 748 1402 800 1411
rect 2554 1402 2606 1454
rect 2640 1402 2692 1454
rect 146 1361 198 1370
rect 146 1327 155 1361
rect 155 1327 189 1361
rect 189 1327 198 1361
rect 146 1318 198 1327
rect 834 1318 886 1370
rect 1350 1361 1402 1370
rect 1350 1327 1359 1361
rect 1359 1327 1393 1361
rect 1393 1327 1402 1361
rect 1350 1318 1402 1327
rect 2038 1361 2090 1370
rect 2038 1327 2047 1361
rect 2047 1327 2081 1361
rect 2081 1327 2090 1361
rect 2038 1318 2090 1327
rect 2554 1361 2606 1370
rect 2554 1327 2563 1361
rect 2563 1327 2597 1361
rect 2597 1327 2606 1361
rect 2554 1318 2606 1327
rect 920 1234 972 1286
rect 1436 1234 1488 1286
rect 748 605 800 614
rect 748 571 757 605
rect 757 571 791 605
rect 791 571 800 605
rect 748 562 800 571
rect 1436 605 1488 614
rect 1436 571 1445 605
rect 1445 571 1479 605
rect 1479 571 1488 605
rect 1436 562 1488 571
rect 2296 562 2348 614
rect 146 142 198 194
rect 920 185 972 194
rect 920 151 929 185
rect 929 151 963 185
rect 963 151 972 185
rect 920 142 972 151
rect 1350 142 1402 194
rect 2038 142 2090 194
rect 2554 142 2606 194
rect 834 58 886 110
rect 920 58 972 110
rect 1264 17 1316 26
rect 1264 -17 1273 17
rect 1273 -17 1307 17
rect 1307 -17 1316 17
rect 1264 -26 1316 -17
rect 2640 17 2692 26
rect 2640 -17 2649 17
rect 2649 -17 2683 17
rect 2683 -17 2692 17
rect 2640 -26 2692 -17
<< metal2 >>
rect 316 2882 372 2888
rect 316 2830 318 2882
rect 370 2830 372 2882
rect 144 1792 200 1801
rect 144 1370 200 1736
rect 316 1792 372 2830
rect 316 1727 372 1736
rect 832 2882 888 2888
rect 832 2830 834 2882
rect 886 2830 888 2882
rect 832 1792 888 2830
rect 1348 2882 1404 2888
rect 1348 2830 1350 2882
rect 1402 2830 1404 2882
rect 832 1727 888 1736
rect 1262 1792 1318 1801
rect 230 1706 286 1712
rect 230 1654 232 1706
rect 284 1654 286 1706
rect 230 1454 286 1654
rect 832 1622 888 1628
rect 832 1570 834 1622
rect 886 1570 888 1622
rect 230 1402 232 1454
rect 284 1402 286 1454
rect 230 1396 286 1402
rect 746 1538 802 1544
rect 746 1486 748 1538
rect 800 1486 802 1538
rect 746 1454 802 1486
rect 746 1402 748 1454
rect 800 1402 802 1454
rect 144 1318 146 1370
rect 198 1318 200 1370
rect 144 194 200 1318
rect 746 614 802 1402
rect 832 1370 888 1570
rect 832 1318 834 1370
rect 886 1318 888 1370
rect 832 1312 888 1318
rect 746 562 748 614
rect 800 562 802 614
rect 746 556 802 562
rect 918 1286 974 1292
rect 918 1234 920 1286
rect 972 1234 974 1286
rect 144 142 146 194
rect 198 142 200 194
rect 144 136 200 142
rect 918 194 974 1234
rect 1262 1288 1318 1736
rect 1348 1790 1404 2830
rect 2036 2882 2092 2888
rect 2036 2830 2038 2882
rect 2090 2830 2092 2882
rect 1348 1738 1350 1790
rect 1402 1738 1404 1790
rect 1348 1706 1404 1738
rect 1348 1654 1350 1706
rect 1402 1654 1404 1706
rect 1348 1648 1404 1654
rect 1434 2462 1490 2468
rect 1434 2410 1436 2462
rect 1488 2410 1490 2462
rect 1262 1223 1318 1232
rect 1348 1370 1404 1376
rect 1348 1318 1350 1370
rect 1402 1318 1404 1370
rect 1348 1288 1404 1318
rect 918 142 920 194
rect 972 142 974 194
rect 832 110 888 116
rect 832 58 834 110
rect 886 58 888 110
rect 832 28 888 58
rect 918 110 974 142
rect 1348 194 1404 1232
rect 1434 1286 1490 2410
rect 2036 1706 2092 2830
rect 2552 2882 2608 2888
rect 2552 2830 2554 2882
rect 2606 2830 2608 2882
rect 2036 1654 2038 1706
rect 2090 1654 2092 1706
rect 2036 1622 2092 1654
rect 2294 2462 2350 2468
rect 2294 2410 2296 2462
rect 2348 2410 2350 2462
rect 2036 1570 2038 1622
rect 2090 1570 2092 1622
rect 2036 1564 2092 1570
rect 2122 1622 2178 1628
rect 2122 1570 2124 1622
rect 2176 1570 2178 1622
rect 1434 1234 1436 1286
rect 1488 1234 1490 1286
rect 1434 614 1490 1234
rect 1434 562 1436 614
rect 1488 562 1490 614
rect 1434 556 1490 562
rect 2036 1370 2092 1376
rect 2036 1318 2038 1370
rect 2090 1318 2092 1370
rect 2036 1288 2092 1318
rect 1348 142 1350 194
rect 1402 142 1404 194
rect 1348 136 1404 142
rect 2036 194 2092 1232
rect 2036 142 2038 194
rect 2090 142 2092 194
rect 2036 136 2092 142
rect 918 58 920 110
rect 972 58 974 110
rect 918 52 974 58
rect 832 -37 888 -28
rect 1262 28 1318 48
rect 1262 -37 1318 -28
rect 2122 28 2178 1570
rect 2294 1538 2350 2410
rect 2552 1706 2608 2830
rect 2552 1654 2554 1706
rect 2606 1654 2608 1706
rect 2552 1622 2608 1654
rect 2552 1570 2554 1622
rect 2606 1570 2608 1622
rect 2552 1564 2608 1570
rect 2638 1792 2694 1801
rect 2294 1486 2296 1538
rect 2348 1486 2350 1538
rect 2294 614 2350 1486
rect 2294 562 2296 614
rect 2348 562 2350 614
rect 2294 556 2350 562
rect 2552 1454 2608 1460
rect 2552 1402 2554 1454
rect 2606 1402 2608 1454
rect 2552 1370 2608 1402
rect 2638 1454 2694 1736
rect 2638 1402 2640 1454
rect 2692 1402 2694 1454
rect 2638 1396 2694 1402
rect 2552 1318 2554 1370
rect 2606 1318 2608 1370
rect 2552 194 2608 1318
rect 2552 142 2554 194
rect 2606 142 2608 194
rect 2552 136 2608 142
rect 2122 -37 2178 -28
rect 2638 28 2694 48
rect 2638 -37 2694 -28
<< via2 >>
rect 144 1736 200 1792
rect 316 1736 372 1792
rect 832 1736 888 1792
rect 1262 1736 1318 1792
rect 1262 1232 1318 1288
rect 1348 1232 1404 1288
rect 2036 1232 2092 1288
rect 832 -28 888 28
rect 1262 26 1318 28
rect 1262 -26 1264 26
rect 1264 -26 1316 26
rect 1316 -26 1318 26
rect 1262 -28 1318 -26
rect 2638 1736 2694 1792
rect 2122 -28 2178 28
rect 2638 26 2694 28
rect 2638 -26 2640 26
rect 2640 -26 2692 26
rect 2692 -26 2694 26
rect 2638 -28 2694 -26
<< metal3 >>
rect -80 1796 2832 1844
rect -80 1792 2040 1796
rect -80 1736 144 1792
rect 200 1736 316 1792
rect 372 1736 832 1792
rect 888 1736 1262 1792
rect 1318 1736 2040 1792
rect -80 1732 2040 1736
rect 2104 1732 2336 1796
rect 2400 1792 2832 1796
rect 2400 1736 2638 1792
rect 2694 1736 2832 1792
rect 2400 1732 2832 1736
rect -80 1684 2832 1732
rect 1257 1288 1409 1340
rect 1257 1232 1262 1288
rect 1318 1232 1348 1288
rect 1404 1232 1409 1288
rect 1257 1180 1409 1232
rect 2031 1292 2105 1340
rect 2031 1288 2040 1292
rect 2031 1232 2036 1288
rect 2031 1228 2040 1232
rect 2104 1228 2105 1292
rect 2031 1180 2105 1228
rect -80 32 2832 80
rect -80 -32 -32 32
rect 32 28 2832 32
rect 32 -28 832 28
rect 888 -28 1262 28
rect 1318 -28 2122 28
rect 2178 -28 2638 28
rect 2694 -28 2832 28
rect 32 -32 2832 -28
rect -80 -80 2832 -32
<< via3 >>
rect 2040 1732 2104 1796
rect 2336 1732 2400 1796
rect 2040 1288 2104 1292
rect 2040 1232 2092 1288
rect 2092 1232 2104 1288
rect 2040 1228 2104 1232
rect -32 -32 32 32
<< metal4 >>
rect -118 32 118 1882
rect 1954 1796 2190 1797
rect 1954 1732 2040 1796
rect 2104 1732 2190 1796
rect 1954 1292 2190 1732
rect 1954 1228 2040 1292
rect 2104 1228 2190 1292
rect 1954 1227 2190 1228
rect 2250 1796 2486 1882
rect 2250 1732 2336 1796
rect 2400 1732 2486 1796
rect -118 -32 -32 32
rect 32 -32 118 32
rect -118 -118 118 -32
rect 2250 -118 2486 1732
<< end >>
