MACRO RING_OSCILLATOR
  ORIGIN 0 0 ;
  FOREIGN RING_OSCILLATOR 0 0 ;
  SIZE 13.02 BY 15.71 ;
  PIN INP
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
      LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
      LAYER M2 ;
        RECT 3.71 2.8 4.03 3.08 ;
      LAYER M3 ;
        RECT 3.73 2.94 4.01 12.18 ;
      LAYER M2 ;
        RECT 3.71 12.04 4.03 12.32 ;
      LAYER M2 ;
        RECT 1.12 7 2.32 7.28 ;
      LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
      LAYER M2 ;
        RECT 1.99 7 2.31 7.28 ;
      LAYER M1 ;
        RECT 2.025 7.14 2.275 7.98 ;
      LAYER M2 ;
        RECT 1.99 7.84 2.31 8.12 ;
      LAYER M3 ;
        RECT 3.73 7.375 4.01 7.745 ;
      LAYER M2 ;
        RECT 2.15 7.42 3.87 7.7 ;
      LAYER M1 ;
        RECT 2.025 7.475 2.275 7.645 ;
    END
  END INP
  OBS 
  LAYER M2 ;
        RECT 1.12 2.8 2.32 3.08 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M2 ;
        RECT 1.13 2.8 1.45 3.08 ;
  LAYER M3 ;
        RECT 1.15 2.94 1.43 12.18 ;
  LAYER M2 ;
        RECT 1.13 12.04 1.45 12.32 ;
  LAYER M2 ;
        RECT 5.42 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 5.42 7.84 6.62 8.12 ;
  LAYER M2 ;
        RECT 5.43 7 5.75 7.28 ;
  LAYER M1 ;
        RECT 5.465 7.14 5.715 7.98 ;
  LAYER M2 ;
        RECT 5.43 7.84 5.75 8.12 ;
  LAYER M3 ;
        RECT 1.15 7.375 1.43 7.745 ;
  LAYER M4 ;
        RECT 1.29 7.16 4.73 7.96 ;
  LAYER M3 ;
        RECT 4.59 7.439 4.87 7.681 ;
  LAYER M2 ;
        RECT 4.73 7.42 5.59 7.7 ;
  LAYER M1 ;
        RECT 5.465 7.475 5.715 7.645 ;
  LAYER M1 ;
        RECT 5.465 7.475 5.715 7.645 ;
  LAYER M2 ;
        RECT 5.42 7.42 5.76 7.7 ;
  LAYER M2 ;
        RECT 4.57 7.42 4.89 7.7 ;
  LAYER M3 ;
        RECT 4.59 7.4 4.87 7.72 ;
  LAYER M3 ;
        RECT 1.15 7.375 1.43 7.745 ;
  LAYER M4 ;
        RECT 1.125 7.16 1.455 7.96 ;
  LAYER M3 ;
        RECT 4.59 7.375 4.87 7.745 ;
  LAYER M4 ;
        RECT 4.565 7.16 4.895 7.96 ;
  LAYER M1 ;
        RECT 5.465 7.475 5.715 7.645 ;
  LAYER M2 ;
        RECT 5.42 7.42 5.76 7.7 ;
  LAYER M3 ;
        RECT 1.15 7.375 1.43 7.745 ;
  LAYER M4 ;
        RECT 1.125 7.16 1.455 7.96 ;
  LAYER M2 ;
        RECT 5.42 2.8 6.62 3.08 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 5.42 12.04 6.62 12.32 ;
  LAYER M2 ;
        RECT 5.43 2.8 5.75 3.08 ;
  LAYER M1 ;
        RECT 5.465 2.94 5.715 6.3 ;
  LAYER M2 ;
        RECT 4.73 6.16 5.59 6.44 ;
  LAYER M1 ;
        RECT 4.605 6.3 4.855 7.14 ;
  LAYER M2 ;
        RECT 4.57 7 4.89 7.28 ;
  LAYER M1 ;
        RECT 4.605 7.14 4.855 7.98 ;
  LAYER M2 ;
        RECT 4.57 7.84 4.89 8.12 ;
  LAYER M1 ;
        RECT 4.605 7.98 4.855 11.76 ;
  LAYER M2 ;
        RECT 4.73 11.62 5.59 11.9 ;
  LAYER M1 ;
        RECT 5.465 11.76 5.715 12.18 ;
  LAYER M2 ;
        RECT 5.43 12.04 5.75 12.32 ;
  LAYER M1 ;
        RECT 4.605 6.215 4.855 6.385 ;
  LAYER M2 ;
        RECT 4.56 6.16 4.9 6.44 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 5.465 2.855 5.715 3.025 ;
  LAYER M2 ;
        RECT 5.42 2.8 5.76 3.08 ;
  LAYER M1 ;
        RECT 5.465 6.215 5.715 6.385 ;
  LAYER M2 ;
        RECT 5.42 6.16 5.76 6.44 ;
  LAYER M1 ;
        RECT 4.605 6.215 4.855 6.385 ;
  LAYER M2 ;
        RECT 4.56 6.16 4.9 6.44 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 5.465 2.855 5.715 3.025 ;
  LAYER M2 ;
        RECT 5.42 2.8 5.76 3.08 ;
  LAYER M1 ;
        RECT 5.465 6.215 5.715 6.385 ;
  LAYER M2 ;
        RECT 5.42 6.16 5.76 6.44 ;
  LAYER M1 ;
        RECT 4.605 6.215 4.855 6.385 ;
  LAYER M2 ;
        RECT 4.56 6.16 4.9 6.44 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.065 ;
  LAYER M2 ;
        RECT 4.56 7.84 4.9 8.12 ;
  LAYER M1 ;
        RECT 5.465 2.855 5.715 3.025 ;
  LAYER M2 ;
        RECT 5.42 2.8 5.76 3.08 ;
  LAYER M1 ;
        RECT 5.465 6.215 5.715 6.385 ;
  LAYER M2 ;
        RECT 5.42 6.16 5.76 6.44 ;
  LAYER M1 ;
        RECT 4.605 6.215 4.855 6.385 ;
  LAYER M2 ;
        RECT 4.56 6.16 4.9 6.44 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.065 ;
  LAYER M2 ;
        RECT 4.56 7.84 4.9 8.12 ;
  LAYER M1 ;
        RECT 5.465 2.855 5.715 3.025 ;
  LAYER M2 ;
        RECT 5.42 2.8 5.76 3.08 ;
  LAYER M1 ;
        RECT 5.465 6.215 5.715 6.385 ;
  LAYER M2 ;
        RECT 5.42 6.16 5.76 6.44 ;
  LAYER M1 ;
        RECT 4.605 6.215 4.855 6.385 ;
  LAYER M2 ;
        RECT 4.56 6.16 4.9 6.44 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.065 ;
  LAYER M2 ;
        RECT 4.56 7.84 4.9 8.12 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 11.845 ;
  LAYER M2 ;
        RECT 4.56 11.62 4.9 11.9 ;
  LAYER M1 ;
        RECT 5.465 2.855 5.715 3.025 ;
  LAYER M2 ;
        RECT 5.42 2.8 5.76 3.08 ;
  LAYER M1 ;
        RECT 5.465 6.215 5.715 6.385 ;
  LAYER M2 ;
        RECT 5.42 6.16 5.76 6.44 ;
  LAYER M1 ;
        RECT 5.465 11.675 5.715 11.845 ;
  LAYER M2 ;
        RECT 5.42 11.62 5.76 11.9 ;
  LAYER M1 ;
        RECT 5.465 12.095 5.715 12.265 ;
  LAYER M2 ;
        RECT 5.42 12.04 5.76 12.32 ;
  LAYER M1 ;
        RECT 4.605 6.215 4.855 6.385 ;
  LAYER M2 ;
        RECT 4.56 6.16 4.9 6.44 ;
  LAYER M1 ;
        RECT 4.605 7.055 4.855 7.225 ;
  LAYER M2 ;
        RECT 4.56 7 4.9 7.28 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.065 ;
  LAYER M2 ;
        RECT 4.56 7.84 4.9 8.12 ;
  LAYER M1 ;
        RECT 4.605 11.675 4.855 11.845 ;
  LAYER M2 ;
        RECT 4.56 11.62 4.9 11.9 ;
  LAYER M1 ;
        RECT 5.465 2.855 5.715 3.025 ;
  LAYER M2 ;
        RECT 5.42 2.8 5.76 3.08 ;
  LAYER M1 ;
        RECT 5.465 6.215 5.715 6.385 ;
  LAYER M2 ;
        RECT 5.42 6.16 5.76 6.44 ;
  LAYER M1 ;
        RECT 5.465 11.675 5.715 11.845 ;
  LAYER M2 ;
        RECT 5.42 11.62 5.76 11.9 ;
  LAYER M1 ;
        RECT 5.465 12.095 5.715 12.265 ;
  LAYER M2 ;
        RECT 5.42 12.04 5.76 12.32 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 5.85 6.58 7.05 6.86 ;
  LAYER M2 ;
        RECT 5.85 0.7 7.05 0.98 ;
  LAYER M2 ;
        RECT 5.42 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 5.42 2.8 6.62 3.08 ;
  LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
  LAYER M1 ;
        RECT 3.745 7.895 3.995 11.425 ;
  LAYER M1 ;
        RECT 3.745 11.675 3.995 12.685 ;
  LAYER M1 ;
        RECT 3.745 13.775 3.995 14.785 ;
  LAYER M1 ;
        RECT 4.175 7.895 4.425 11.425 ;
  LAYER M1 ;
        RECT 3.315 7.895 3.565 11.425 ;
  LAYER M2 ;
        RECT 3.27 8.26 4.47 8.54 ;
  LAYER M2 ;
        RECT 3.27 14.14 4.47 14.42 ;
  LAYER M2 ;
        RECT 3.7 7.84 4.9 8.12 ;
  LAYER M2 ;
        RECT 3.7 12.04 4.9 12.32 ;
  LAYER M3 ;
        RECT 3.3 8.24 3.58 14.44 ;
  LAYER M1 ;
        RECT 6.325 7.895 6.575 11.425 ;
  LAYER M1 ;
        RECT 6.325 11.675 6.575 12.685 ;
  LAYER M1 ;
        RECT 6.325 13.775 6.575 14.785 ;
  LAYER M1 ;
        RECT 5.895 7.895 6.145 11.425 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M2 ;
        RECT 5.85 8.26 7.05 8.54 ;
  LAYER M2 ;
        RECT 5.85 14.14 7.05 14.42 ;
  LAYER M2 ;
        RECT 5.42 7.84 6.62 8.12 ;
  LAYER M2 ;
        RECT 5.42 12.04 6.62 12.32 ;
  LAYER M3 ;
        RECT 6.74 8.24 7.02 14.44 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 1.12 7 2.32 7.28 ;
  LAYER M2 ;
        RECT 1.12 2.8 2.32 3.08 ;
  LAYER M3 ;
        RECT 0.72 0.68 1 6.88 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 1.12 7.84 2.32 8.12 ;
  LAYER M2 ;
        RECT 1.12 12.04 2.32 12.32 ;
  LAYER M3 ;
        RECT 0.72 8.24 1 14.44 ;
  END 
END RING_OSCILLATOR
