magic
tech sky130A
magscale 1 2
timestamp 1677423745
<< locali >>
rect 405 1579 413 1613
rect 447 1579 455 1613
rect 405 1445 455 1579
rect 405 1411 413 1445
rect 447 1411 455 1445
<< viali >>
rect 413 1579 447 1613
rect 413 1411 447 1445
<< metal1 >>
rect 226 2462 290 2464
rect 226 2410 232 2462
rect 284 2410 290 2462
rect 226 2408 290 2410
rect 396 1613 464 1624
rect 396 1579 413 1613
rect 447 1579 464 1613
rect 396 1568 464 1579
rect 396 1445 464 1456
rect 396 1411 413 1445
rect 447 1411 464 1445
rect 396 1400 464 1411
rect 226 614 290 616
rect 226 562 232 614
rect 284 562 290 614
rect 226 560 290 562
<< via1 >>
rect 232 2410 284 2462
rect 232 562 284 614
<< metal2 >>
rect 230 2462 286 2468
rect 230 2410 232 2462
rect 284 2410 286 2462
rect 230 614 286 2410
rect 230 562 232 614
rect 284 562 286 614
rect 230 556 286 562
use NMOS_S_25628869_X1_Y1_1677407590_1677407590  NMOS_S_25628869_X1_Y1_1677407590_1677407590_0
timestamp 1677423745
transform -1 0 516 0 -1 1512
box 52 56 395 1482
use PMOS_S_89421238_X1_Y1_1677407591_1677407590  PMOS_S_89421238_X1_Y1_1677407591_1677407590_0
timestamp 1677423745
transform -1 0 516 0 1 1512
box 0 0 516 1512
<< end >>
