MACRO ANALOG
  ORIGIN 0 0 ;
  FOREIGN ANALOG 0 0 ;
  SIZE 13.02 BY 23.27 ;
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M4 ;
        RECT 3.275 5.9 5.325 6.7 ;
      LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
      LAYER M2 ;
        RECT 6.28 7.84 7.48 8.12 ;
      LAYER M2 ;
        RECT 6.29 7 6.61 7.28 ;
      LAYER M1 ;
        RECT 6.325 7.14 6.575 7.98 ;
      LAYER M2 ;
        RECT 6.29 7.84 6.61 8.12 ;
      LAYER M2 ;
        RECT 3.7 10.36 4.9 10.64 ;
      LAYER M2 ;
        RECT 1.98 10.36 3.18 10.64 ;
      LAYER M4 ;
        RECT 4.995 5.9 5.325 6.7 ;
      LAYER M3 ;
        RECT 5.02 6.3 5.3 7.14 ;
      LAYER M2 ;
        RECT 5.16 7 6.45 7.28 ;
      LAYER M2 ;
        RECT 5 7 5.32 7.28 ;
      LAYER M1 ;
        RECT 5.035 7.14 5.285 10.5 ;
      LAYER M2 ;
        RECT 4.73 10.36 5.16 10.64 ;
      LAYER M2 ;
        RECT 3.01 10.36 3.87 10.64 ;
    END
  END Y
  OBS 
  LAYER M4 ;
        RECT 0.695 4.64 2.745 5.44 ;
  LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
  LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
  LAYER M2 ;
        RECT 6.29 2.8 6.61 3.08 ;
  LAYER M3 ;
        RECT 6.31 2.94 6.59 12.18 ;
  LAYER M2 ;
        RECT 6.29 12.04 6.61 12.32 ;
  LAYER M2 ;
        RECT 1.12 15.4 2.32 15.68 ;
  LAYER M2 ;
        RECT 5.85 15.4 7.05 15.68 ;
  LAYER M4 ;
        RECT 2.58 4.64 3.44 5.44 ;
  LAYER M3 ;
        RECT 3.3 4.919 3.58 5.161 ;
  LAYER M2 ;
        RECT 3.44 4.9 6.45 5.18 ;
  LAYER M3 ;
        RECT 6.31 4.855 6.59 5.225 ;
  LAYER M2 ;
        RECT 3.01 12.04 6.45 12.32 ;
  LAYER M1 ;
        RECT 2.885 12.18 3.135 15.54 ;
  LAYER M2 ;
        RECT 2.15 15.4 3.01 15.68 ;
  LAYER M2 ;
        RECT 3.01 15.4 6.02 15.68 ;
  LAYER M2 ;
        RECT 3.28 4.9 3.6 5.18 ;
  LAYER M3 ;
        RECT 3.3 4.88 3.58 5.2 ;
  LAYER M2 ;
        RECT 6.29 4.9 6.61 5.18 ;
  LAYER M3 ;
        RECT 6.31 4.88 6.59 5.2 ;
  LAYER M3 ;
        RECT 3.3 4.855 3.58 5.225 ;
  LAYER M4 ;
        RECT 3.275 4.64 3.605 5.44 ;
  LAYER M2 ;
        RECT 6.29 4.9 6.61 5.18 ;
  LAYER M3 ;
        RECT 6.31 4.88 6.59 5.2 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 12.265 ;
  LAYER M2 ;
        RECT 2.84 12.04 3.18 12.32 ;
  LAYER M1 ;
        RECT 2.885 15.455 3.135 15.625 ;
  LAYER M2 ;
        RECT 2.84 15.4 3.18 15.68 ;
  LAYER M2 ;
        RECT 6.29 4.9 6.61 5.18 ;
  LAYER M3 ;
        RECT 6.31 4.88 6.59 5.2 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 12.265 ;
  LAYER M2 ;
        RECT 2.84 12.04 3.18 12.32 ;
  LAYER M1 ;
        RECT 2.885 15.455 3.135 15.625 ;
  LAYER M2 ;
        RECT 2.84 15.4 3.18 15.68 ;
  LAYER M2 ;
        RECT 6.29 4.9 6.61 5.18 ;
  LAYER M3 ;
        RECT 6.31 4.88 6.59 5.2 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 12.265 ;
  LAYER M2 ;
        RECT 2.84 12.04 3.18 12.32 ;
  LAYER M1 ;
        RECT 2.885 15.455 3.135 15.625 ;
  LAYER M2 ;
        RECT 2.84 15.4 3.18 15.68 ;
  LAYER M2 ;
        RECT 6.29 4.9 6.61 5.18 ;
  LAYER M3 ;
        RECT 6.31 4.88 6.59 5.2 ;
  LAYER M1 ;
        RECT 2.885 12.095 3.135 12.265 ;
  LAYER M2 ;
        RECT 2.84 12.04 3.18 12.32 ;
  LAYER M1 ;
        RECT 2.885 15.455 3.135 15.625 ;
  LAYER M2 ;
        RECT 2.84 15.4 3.18 15.68 ;
  LAYER M2 ;
        RECT 6.29 4.9 6.61 5.18 ;
  LAYER M3 ;
        RECT 6.31 4.88 6.59 5.2 ;
  LAYER M2 ;
        RECT 1.98 14.56 3.18 14.84 ;
  LAYER M2 ;
        RECT 3.7 14.56 4.9 14.84 ;
  LAYER M4 ;
        RECT 2.845 15.98 4.895 16.78 ;
  LAYER M2 ;
        RECT 1.12 19.6 2.32 19.88 ;
  LAYER M2 ;
        RECT 5.85 19.6 7.05 19.88 ;
  LAYER M2 ;
        RECT 3.01 14.56 3.87 14.84 ;
  LAYER M2 ;
        RECT 2.85 14.56 3.17 14.84 ;
  LAYER M3 ;
        RECT 2.87 14.7 3.15 16.38 ;
  LAYER M4 ;
        RECT 2.845 15.98 3.175 16.78 ;
  LAYER M3 ;
        RECT 2.87 16.38 3.15 19.74 ;
  LAYER M2 ;
        RECT 2.15 19.6 3.01 19.88 ;
  LAYER M2 ;
        RECT 3.01 19.6 6.02 19.88 ;
  LAYER M2 ;
        RECT 2.85 14.56 3.17 14.84 ;
  LAYER M3 ;
        RECT 2.87 14.54 3.15 14.86 ;
  LAYER M3 ;
        RECT 2.87 16.195 3.15 16.565 ;
  LAYER M4 ;
        RECT 2.845 15.98 3.175 16.78 ;
  LAYER M2 ;
        RECT 2.85 14.56 3.17 14.84 ;
  LAYER M3 ;
        RECT 2.87 14.54 3.15 14.86 ;
  LAYER M3 ;
        RECT 2.87 16.195 3.15 16.565 ;
  LAYER M4 ;
        RECT 2.845 15.98 3.175 16.78 ;
  LAYER M2 ;
        RECT 2.85 14.56 3.17 14.84 ;
  LAYER M3 ;
        RECT 2.87 14.54 3.15 14.86 ;
  LAYER M2 ;
        RECT 2.85 19.6 3.17 19.88 ;
  LAYER M3 ;
        RECT 2.87 19.58 3.15 19.9 ;
  LAYER M3 ;
        RECT 2.87 16.195 3.15 16.565 ;
  LAYER M4 ;
        RECT 2.845 15.98 3.175 16.78 ;
  LAYER M2 ;
        RECT 2.85 14.56 3.17 14.84 ;
  LAYER M3 ;
        RECT 2.87 14.54 3.15 14.86 ;
  LAYER M2 ;
        RECT 2.85 19.6 3.17 19.88 ;
  LAYER M3 ;
        RECT 2.87 19.58 3.15 19.9 ;
  LAYER M3 ;
        RECT 2.87 16.195 3.15 16.565 ;
  LAYER M4 ;
        RECT 2.845 15.98 3.175 16.78 ;
  LAYER M2 ;
        RECT 2.85 14.56 3.17 14.84 ;
  LAYER M3 ;
        RECT 2.87 14.54 3.15 14.86 ;
  LAYER M2 ;
        RECT 2.85 19.6 3.17 19.88 ;
  LAYER M3 ;
        RECT 2.87 19.58 3.15 19.9 ;
  LAYER M3 ;
        RECT 2.87 16.195 3.15 16.565 ;
  LAYER M4 ;
        RECT 2.845 15.98 3.175 16.78 ;
  LAYER M2 ;
        RECT 2.85 14.56 3.17 14.84 ;
  LAYER M3 ;
        RECT 2.87 14.54 3.15 14.86 ;
  LAYER M2 ;
        RECT 2.85 19.6 3.17 19.88 ;
  LAYER M3 ;
        RECT 2.87 19.58 3.15 19.9 ;
  LAYER M3 ;
        RECT 2.87 16.195 3.15 16.565 ;
  LAYER M4 ;
        RECT 2.845 15.98 3.175 16.78 ;
  LAYER M1 ;
        RECT 7.185 3.695 7.435 7.225 ;
  LAYER M1 ;
        RECT 7.185 2.435 7.435 3.445 ;
  LAYER M1 ;
        RECT 7.185 0.335 7.435 1.345 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M1 ;
        RECT 7.615 3.695 7.865 7.225 ;
  LAYER M2 ;
        RECT 6.71 0.7 7.91 0.98 ;
  LAYER M2 ;
        RECT 6.71 6.58 7.91 6.86 ;
  LAYER M2 ;
        RECT 6.28 7 7.48 7.28 ;
  LAYER M2 ;
        RECT 6.28 2.8 7.48 3.08 ;
  LAYER M3 ;
        RECT 7.6 0.68 7.88 6.88 ;
  LAYER M1 ;
        RECT 7.185 7.895 7.435 11.425 ;
  LAYER M1 ;
        RECT 7.185 11.675 7.435 12.685 ;
  LAYER M1 ;
        RECT 7.185 13.775 7.435 14.785 ;
  LAYER M1 ;
        RECT 6.755 7.895 7.005 11.425 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M2 ;
        RECT 6.71 14.14 7.91 14.42 ;
  LAYER M2 ;
        RECT 6.71 8.26 7.91 8.54 ;
  LAYER M2 ;
        RECT 6.28 7.84 7.48 8.12 ;
  LAYER M2 ;
        RECT 6.28 12.04 7.48 12.32 ;
  LAYER M3 ;
        RECT 7.6 8.24 7.88 14.44 ;
  LAYER M4 ;
        RECT 3.44 17.75 4.74 19.05 ;
  LAYER M4 ;
        RECT 4.29 16.58 4.74 19.1 ;
  LAYER M5 ;
        RECT 3.665 18.07 4.115 20.59 ;
  LAYER M4 ;
        RECT 2.845 19.76 4.895 20.56 ;
  LAYER M4 ;
        RECT 2.845 15.98 4.895 16.78 ;
  LAYER M4 ;
        RECT 0.85 2.37 2.15 3.67 ;
  LAYER M4 ;
        RECT 0.85 2.32 1.3 4.84 ;
  LAYER M5 ;
        RECT 1.475 0.83 1.925 3.35 ;
  LAYER M4 ;
        RECT 0.695 0.86 2.745 1.66 ;
  LAYER M4 ;
        RECT 0.695 4.64 2.745 5.44 ;
  LAYER M4 ;
        RECT 3.87 3.63 5.17 4.93 ;
  LAYER M4 ;
        RECT 4.72 3.58 5.17 6.1 ;
  LAYER M5 ;
        RECT 4.095 2.09 4.545 4.61 ;
  LAYER M4 ;
        RECT 3.275 2.12 5.325 2.92 ;
  LAYER M4 ;
        RECT 3.275 5.9 5.325 6.7 ;
  LAYER M1 ;
        RECT 2.025 11.255 2.275 14.785 ;
  LAYER M1 ;
        RECT 2.025 9.995 2.275 11.005 ;
  LAYER M1 ;
        RECT 2.025 7.895 2.275 8.905 ;
  LAYER M1 ;
        RECT 2.455 11.255 2.705 14.785 ;
  LAYER M1 ;
        RECT 1.595 11.255 1.845 14.785 ;
  LAYER M2 ;
        RECT 1.55 8.26 2.75 8.54 ;
  LAYER M2 ;
        RECT 1.55 14.14 2.75 14.42 ;
  LAYER M2 ;
        RECT 1.98 14.56 3.18 14.84 ;
  LAYER M2 ;
        RECT 1.98 10.36 3.18 10.64 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M1 ;
        RECT 1.165 15.455 1.415 18.985 ;
  LAYER M1 ;
        RECT 1.165 19.235 1.415 20.245 ;
  LAYER M1 ;
        RECT 1.165 21.335 1.415 22.345 ;
  LAYER M1 ;
        RECT 1.595 15.455 1.845 18.985 ;
  LAYER M1 ;
        RECT 0.735 15.455 0.985 18.985 ;
  LAYER M2 ;
        RECT 0.69 21.7 1.89 21.98 ;
  LAYER M2 ;
        RECT 0.69 15.82 1.89 16.1 ;
  LAYER M2 ;
        RECT 1.12 15.4 2.32 15.68 ;
  LAYER M2 ;
        RECT 1.12 19.6 2.32 19.88 ;
  LAYER M3 ;
        RECT 0.72 15.8 1 22 ;
  LAYER M1 ;
        RECT 6.755 15.455 7.005 18.985 ;
  LAYER M1 ;
        RECT 6.755 19.235 7.005 20.245 ;
  LAYER M1 ;
        RECT 6.755 21.335 7.005 22.345 ;
  LAYER M1 ;
        RECT 6.325 15.455 6.575 18.985 ;
  LAYER M1 ;
        RECT 7.185 15.455 7.435 18.985 ;
  LAYER M2 ;
        RECT 6.28 21.7 7.48 21.98 ;
  LAYER M2 ;
        RECT 6.28 15.82 7.48 16.1 ;
  LAYER M2 ;
        RECT 5.85 15.4 7.05 15.68 ;
  LAYER M2 ;
        RECT 5.85 19.6 7.05 19.88 ;
  LAYER M3 ;
        RECT 7.17 15.8 7.45 22 ;
  LAYER M1 ;
        RECT 4.605 11.255 4.855 14.785 ;
  LAYER M1 ;
        RECT 4.605 9.995 4.855 11.005 ;
  LAYER M1 ;
        RECT 4.605 7.895 4.855 8.905 ;
  LAYER M1 ;
        RECT 4.175 11.255 4.425 14.785 ;
  LAYER M1 ;
        RECT 5.035 11.255 5.285 14.785 ;
  LAYER M2 ;
        RECT 4.13 8.26 5.33 8.54 ;
  LAYER M2 ;
        RECT 4.13 14.14 5.33 14.42 ;
  LAYER M2 ;
        RECT 3.7 14.56 4.9 14.84 ;
  LAYER M2 ;
        RECT 3.7 10.36 4.9 10.64 ;
  LAYER M3 ;
        RECT 5.02 8.24 5.3 14.44 ;
  END 
END ANALOG
