magic
tech sky130A
magscale 1 2
timestamp 1676388708
<< pwell >>
rect 215 1206 301 1482
rect 121 499 395 635
<< nmos >>
rect 200 525 230 609
rect 286 525 316 609
<< ndiff >>
rect 147 575 200 609
rect 147 541 155 575
rect 189 541 200 575
rect 147 525 200 541
rect 230 575 286 609
rect 230 541 241 575
rect 275 541 286 575
rect 230 525 286 541
rect 316 575 369 609
rect 316 541 327 575
rect 361 541 369 575
rect 316 525 369 541
<< ndiffc >>
rect 155 541 189 575
rect 241 541 275 575
rect 327 541 361 575
<< psubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
<< psubdiffcont >>
rect 241 1327 275 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 609 230 897
rect 286 609 316 897
rect 200 252 230 525
rect 286 252 316 525
<< polycont >>
rect 241 907 275 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 147 575 197 773
rect 147 541 155 575
rect 189 541 197 575
rect 147 185 197 541
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 575 283 773
rect 233 541 241 575
rect 275 541 283 575
rect 233 101 283 541
rect 233 67 241 101
rect 275 67 283 101
rect 319 575 369 773
rect 319 541 327 575
rect 361 541 369 575
rect 319 185 369 541
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
<< viali >>
rect 241 1327 275 1361
rect 241 907 275 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
<< metal1 >>
rect 138 1370 378 1372
rect 138 1361 318 1370
rect 138 1327 241 1361
rect 275 1327 318 1361
rect 138 1318 318 1327
rect 370 1318 378 1370
rect 138 1316 378 1318
rect 52 941 292 952
rect 52 907 241 941
rect 275 907 292 941
rect 52 896 292 907
rect 138 194 378 196
rect 138 185 318 194
rect 138 151 155 185
rect 189 151 318 185
rect 138 142 318 151
rect 370 142 378 194
rect 138 140 378 142
rect 52 101 292 112
rect 52 67 241 101
rect 275 67 292 101
rect 52 56 292 67
<< via1 >>
rect 318 1318 370 1370
rect 318 185 370 194
rect 318 151 327 185
rect 327 151 361 185
rect 361 151 370 185
rect 318 142 370 151
<< metal2 >>
rect 316 1370 372 1376
rect 316 1318 318 1370
rect 370 1318 372 1370
rect 316 194 372 1318
rect 316 142 318 194
rect 370 142 372 194
rect 316 136 372 142
<< end >>
