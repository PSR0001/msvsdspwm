* NGSPICE file created from TEST_0.ext - technology: sky130A

.subckt PMOS_S_95137167_X1_Y1_1676553145_1676553145 a_200_252# a_230_399# w_0_0#
X0 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=3.92e+06u as=8.904e+11p ps=7.78e+06u w=1.68e+06u l=150000u
X1 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
C0 a_230_399# w_0_0# 0.78fF
C1 w_0_0# a_200_252# 0.66fF
C2 a_230_399# a_200_252# 0.10fF
C3 a_230_399# VSUBS -0.03fF
C4 a_200_252# VSUBS 0.06fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt NMOS_S_54129001_X1_Y1_1676553144_1676553145 a_200_252# a_230_483# a_147_483#
X0 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_200_252# a_230_483# 0.11fF
C1 a_230_483# a_147_483# 0.74fF
C2 a_200_252# a_147_483# 0.89fF
.ends

.subckt INV_45746474_0_0_1676553145 PMOS_S_95137167_X1_Y1_1676553145_1676553145_0/w_0_0#
+ m1_398_560# li_405_1411# VSUBS
XPMOS_S_95137167_X1_Y1_1676553145_1676553145_0 m1_398_560# li_405_1411# PMOS_S_95137167_X1_Y1_1676553145_1676553145_0/w_0_0#
+ PMOS_S_95137167_X1_Y1_1676553145_1676553145
XNMOS_S_54129001_X1_Y1_1676553144_1676553145_0 m1_398_560# li_405_1411# VSUBS NMOS_S_54129001_X1_Y1_1676553144_1676553145
C0 li_405_1411# PMOS_S_95137167_X1_Y1_1676553145_1676553145_0/w_0_0# 0.06fF
C1 PMOS_S_95137167_X1_Y1_1676553145_1676553145_0/w_0_0# m1_398_560# 0.28fF
C2 li_405_1411# m1_398_560# 0.15fF
C3 li_405_1411# VSUBS 0.69fF
C4 m1_398_560# VSUBS 1.53fF
C5 PMOS_S_95137167_X1_Y1_1676553145_1676553145_0/w_0_0# VSUBS 3.02fF
.ends

.subckt DP_PMOS_83764739_X1_Y1_1676553146 a_372_252# a_200_252# a_230_399# a_402_399#
+ w_0_0#
X0 w_0_0# a_372_252# a_402_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=1.3608e+12p pd=1.17e+07u as=4.704e+11p ps=3.92e+06u w=1.68e+06u l=150000u
X1 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=3.92e+06u as=0p ps=0u w=1.68e+06u l=150000u
X2 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
X3 a_402_399# a_372_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
C0 a_200_252# a_230_399# 0.10fF
C1 a_230_399# w_0_0# 0.72fF
C2 a_200_252# a_402_399# 0.01fF
C3 a_372_252# a_402_399# 0.10fF
C4 a_402_399# w_0_0# 0.91fF
C5 a_200_252# a_372_252# 0.21fF
C6 a_230_399# a_402_399# 0.06fF
C7 a_200_252# w_0_0# 0.56fF
C8 a_372_252# w_0_0# 0.57fF
C9 a_402_399# VSUBS -0.05fF
C10 a_230_399# VSUBS -0.10fF
C11 a_372_252# VSUBS 0.04fF
C12 a_200_252# VSUBS -0.00fF
C13 w_0_0# VSUBS 3.45fF
.ends

.subckt NMOS_S_54129001_X1_Y1_1676553147 a_200_252# a_230_483# a_147_483#
X0 a_230_483# a_200_252# a_147_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=2.352e+11p pd=2.24e+06u as=4.452e+11p ps=4.42e+06u w=840000u l=150000u
X1 a_147_483# a_200_252# a_230_483# a_147_483# sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=840000u l=150000u
C0 a_230_483# a_200_252# 0.11fF
C1 a_230_483# a_147_483# 0.74fF
C2 a_200_252# a_147_483# 0.89fF
.ends

.subckt PMOS_S_95137167_X1_Y1_1676553148 a_200_252# a_230_399# w_0_0#
X0 a_230_399# a_200_252# w_0_0# w_0_0# sky130_fd_pr__pfet_01v8 ad=4.704e+11p pd=3.92e+06u as=8.904e+11p ps=7.78e+06u w=1.68e+06u l=150000u
X1 w_0_0# a_200_252# a_230_399# w_0_0# sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.68e+06u l=150000u
C0 a_200_252# a_230_399# 0.10fF
C1 a_200_252# w_0_0# 0.66fF
C2 a_230_399# w_0_0# 0.78fF
C3 a_230_399# VSUBS -0.03fF
C4 a_200_252# VSUBS 0.06fF
C5 w_0_0# VSUBS 2.97fF
.ends

.subckt TEST_0 F E D C B A VDD VSS Y
XINV_45746474_0_0_1676553145_0 m1_312_224# E Y VSS INV_45746474_0_0_1676553145
XDP_PMOS_83764739_X1_Y1_1676553146_0 li_2813_487# m1_1978_560# VDD VDD VDD DP_PMOS_83764739_X1_Y1_1676553146
XNMOS_S_54129001_X1_Y1_1676553147_0 m1_1806_2408# Y VSS NMOS_S_54129001_X1_Y1_1676553147
XPMOS_S_95137167_X1_Y1_1676553148_0 m1_2838_2408# m1_312_224# VDD PMOS_S_95137167_X1_Y1_1676553148
XNMOS_S_54129001_X1_Y1_1676553147_1 m1_1978_560# Y VSS NMOS_S_54129001_X1_Y1_1676553147
XPMOS_S_95137167_X1_Y1_1676553148_1 C m1_312_224# VDD PMOS_S_95137167_X1_Y1_1676553148
XNMOS_S_54129001_X1_Y1_1676553147_2 F VSS VSS NMOS_S_54129001_X1_Y1_1676553147
XNMOS_S_54129001_X1_Y1_1676553147_3 D VSS VSS NMOS_S_54129001_X1_Y1_1676553147
XPMOS_S_95137167_X1_Y1_1676553148_2 m1_946_560# Y m1_312_224# PMOS_S_95137167_X1_Y1_1676553148
XNMOS_S_54129001_X1_Y1_1676553147_4 B VSS VSS NMOS_S_54129001_X1_Y1_1676553147
C0 E F 0.03fF
C1 li_2813_487# m1_312_224# 0.00fF
C2 B m1_312_224# 0.00fF
C3 Y C 0.00fF
C4 Y m1_1806_2408# 0.00fF
C5 Y F 0.01fF
C6 D B 0.00fF
C7 Y A 0.01fF
C8 m1_2838_2408# m1_1806_2408# 0.00fF
C9 D m1_312_224# 0.00fF
C10 B F 0.00fF
C11 m1_312_224# C 0.01fF
C12 B A 0.00fF
C13 m1_312_224# m1_1806_2408# 0.00fF
C14 F m1_312_224# 0.26fF
C15 m1_312_224# A 0.00fF
C16 D C 0.03fF
C17 m1_1978_560# m1_946_560# 0.00fF
C18 Y VDD 0.07fF
C19 A C 0.00fF
C20 F A 0.03fF
C21 Y m1_946_560# 0.00fF
C22 li_2813_487# VDD 0.01fF
C23 B VDD 0.26fF
C24 VDD m1_312_224# 1.60fF
C25 m1_312_224# m1_946_560# 0.00fF
C26 D VDD 0.15fF
C27 VDD C 0.24fF
C28 F VDD 0.00fF
C29 VDD A 0.18fF
C30 E Y 0.04fF
C31 li_2813_487# m1_1978_560# 0.00fF
C32 E m1_312_224# 0.04fF
C33 m1_1978_560# m1_312_224# 0.00fF
C34 E C 0.01fF
C35 Y m1_312_224# 0.65fF
C37 B VSS 0.46fF
C38 m1_946_560# VSS 0.14fF
C39 D VSS 0.56fF
C40 F VSS 0.38fF
C41 C VSS -0.44fF
C42 m1_2838_2408# VSS 0.15fF
C43 m1_1806_2408# VSS 0.97fF
C44 VDD VSS 9.73fF
C45 li_2813_487# VSS 0.28fF
C46 m1_1978_560# VSS 0.98fF
C47 Y VSS 2.89fF
C48 E VSS 1.17fF
C49 m1_312_224# VSS 4.53fF
.ends
