magic
tech sky130A
magscale 1 2
timestamp 1678383033
<< locali >>
rect 61 1747 69 1781
rect 103 1747 111 1781
rect 61 17 111 1747
rect 577 1747 585 1781
rect 619 1747 627 1781
rect 405 1495 413 1529
rect 447 1495 455 1529
rect 61 -17 69 17
rect 103 -17 111 17
rect 577 17 627 1747
rect 1093 1495 1101 1529
rect 1135 1495 1143 1529
rect 577 -17 585 17
rect 619 -17 627 17
<< viali >>
rect 69 1747 103 1781
rect 585 1747 619 1781
rect 413 1495 447 1529
rect 69 -17 103 17
rect 1101 1495 1135 1529
rect 585 -17 619 17
<< metal1 >>
rect 52 1790 204 1792
rect 52 1781 146 1790
rect 52 1747 69 1781
rect 103 1747 146 1781
rect 52 1738 146 1747
rect 198 1738 204 1790
rect 52 1736 204 1738
rect 568 1790 720 1792
rect 568 1781 662 1790
rect 568 1747 585 1781
rect 619 1747 662 1781
rect 568 1738 662 1747
rect 714 1738 720 1790
rect 568 1736 720 1738
rect 1172 1790 1408 1792
rect 1172 1738 1178 1790
rect 1230 1738 1350 1790
rect 1402 1738 1408 1790
rect 1172 1736 1408 1738
rect 396 1538 806 1540
rect 396 1529 748 1538
rect 396 1495 413 1529
rect 447 1495 748 1529
rect 396 1486 748 1495
rect 800 1486 806 1538
rect 396 1484 806 1486
rect 914 1538 1152 1540
rect 914 1486 920 1538
rect 972 1529 1152 1538
rect 972 1495 1101 1529
rect 1135 1495 1152 1529
rect 972 1486 1152 1495
rect 914 1484 1152 1486
rect 54 1286 204 1288
rect 54 1234 60 1286
rect 112 1234 146 1286
rect 198 1234 204 1286
rect 54 1232 204 1234
rect 570 1286 720 1288
rect 570 1234 576 1286
rect 628 1234 662 1286
rect 714 1234 720 1286
rect 570 1232 720 1234
rect 1258 1286 1408 1288
rect 1258 1234 1264 1286
rect 1316 1234 1350 1286
rect 1402 1234 1408 1286
rect 1258 1232 1408 1234
rect 52 26 120 28
rect 52 -26 60 26
rect 112 -26 120 26
rect 52 -28 120 -26
rect 568 26 636 28
rect 568 -26 576 26
rect 628 -26 636 26
rect 568 -28 636 -26
<< via1 >>
rect 146 1738 198 1790
rect 662 1738 714 1790
rect 1178 1738 1230 1790
rect 1350 1738 1402 1790
rect 748 1486 800 1538
rect 920 1486 972 1538
rect 60 1234 112 1286
rect 146 1234 198 1286
rect 576 1234 628 1286
rect 662 1234 714 1286
rect 1264 1234 1316 1286
rect 1350 1234 1402 1286
rect 60 17 112 26
rect 60 -17 69 17
rect 69 -17 103 17
rect 103 -17 112 17
rect 60 -26 112 -17
rect 576 17 628 26
rect 576 -17 585 17
rect 585 -17 619 17
rect 619 -17 628 17
rect 576 -26 628 -17
<< metal2 >>
rect 58 1792 114 1801
rect 58 1286 114 1736
rect 144 1790 200 1796
rect 144 1738 146 1790
rect 198 1738 200 1790
rect 144 1732 200 1738
rect 574 1792 630 1801
rect 230 1540 286 1549
rect 230 1475 286 1484
rect 58 1234 60 1286
rect 112 1234 114 1286
rect 58 1228 114 1234
rect 144 1286 200 1292
rect 144 1234 146 1286
rect 198 1234 200 1286
rect 144 1228 200 1234
rect 574 1286 630 1736
rect 660 1790 716 1796
rect 660 1738 662 1790
rect 714 1738 716 1790
rect 660 1732 716 1738
rect 1176 1790 1232 1796
rect 1176 1738 1178 1790
rect 1230 1738 1232 1790
rect 746 1538 802 1544
rect 746 1486 748 1538
rect 800 1486 802 1538
rect 746 1480 802 1486
rect 918 1540 974 1549
rect 918 1475 974 1484
rect 574 1234 576 1286
rect 628 1234 630 1286
rect 574 1228 630 1234
rect 660 1286 716 1292
rect 660 1234 662 1286
rect 714 1234 716 1286
rect 660 1228 716 1234
rect 58 28 114 48
rect 58 -37 114 -28
rect 574 28 630 48
rect 574 -37 630 -28
rect 1176 28 1232 1738
rect 1262 1792 1318 1801
rect 1262 1286 1318 1736
rect 1348 1790 1404 1796
rect 1348 1738 1350 1790
rect 1402 1738 1404 1790
rect 1348 1732 1404 1738
rect 1262 1234 1264 1286
rect 1316 1234 1318 1286
rect 1262 1228 1318 1234
rect 1348 1286 1404 1292
rect 1348 1234 1350 1286
rect 1402 1234 1404 1286
rect 1348 1228 1404 1234
rect 1176 -37 1232 -28
<< via2 >>
rect 58 1736 114 1792
rect 574 1736 630 1792
rect 230 1484 286 1540
rect 918 1538 974 1540
rect 918 1486 920 1538
rect 920 1486 972 1538
rect 972 1486 974 1538
rect 918 1484 974 1486
rect 58 26 114 28
rect 58 -26 60 26
rect 60 -26 112 26
rect 112 -26 114 26
rect 58 -28 114 -26
rect 574 26 630 28
rect 574 -26 576 26
rect 576 -26 628 26
rect 628 -26 630 26
rect 574 -28 630 -26
rect 1262 1736 1318 1792
rect 1176 -28 1232 28
<< metal3 >>
rect -80 1796 2448 1844
rect -80 1792 2336 1796
rect -80 1736 58 1792
rect 114 1736 574 1792
rect 630 1736 1262 1792
rect 1318 1736 2336 1792
rect -80 1732 2336 1736
rect 2400 1732 2448 1796
rect -80 1684 2448 1732
rect 225 1540 979 1592
rect 225 1484 230 1540
rect 286 1484 918 1540
rect 974 1484 979 1540
rect 225 1432 979 1484
rect -80 32 2448 80
rect -80 -32 -32 32
rect 32 28 2448 32
rect 32 -28 58 28
rect 114 -28 574 28
rect 630 -28 1176 28
rect 1232 -28 2448 28
rect 32 -32 2448 -28
rect -80 -80 2448 -32
<< via3 >>
rect 2336 1732 2400 1796
rect -32 -32 32 32
<< metal4 >>
rect -118 32 118 1882
rect -118 -32 -32 32
rect 32 -32 118 32
rect -118 -118 118 -32
rect 2250 1796 2486 1882
rect 2250 1732 2336 1796
rect 2400 1732 2486 1796
rect 2250 -118 2486 1732
use INV_49597392_PG0_0_0_1678382967  INV_49597392_PG0_0_0_1678382967_0
timestamp 1678383033
transform -1 0 516 0 1 0
box 0 30 516 3024
use STAGE2_INV_2455088_PG0_0_0_1678382968  STAGE2_INV_2455088_PG0_0_0_1678382968_0
timestamp 1678383033
transform -1 0 1548 0 1 0
box 0 30 1032 3024
<< labels >>
flabel metal1 s 860 588 860 588 0 FreeSerif 0 0 0 0 INP
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal1 s 645 1260 645 1260 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 2368 882 2368 882 0 FreeSerif 0 0 0 0 GND
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal1 s 645 1764 645 1764 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
flabel metal4 s 0 882 0 882 0 FreeSerif 0 0 0 0 VCC
<< end >>
