magic
tech sky130A
magscale 1 2
timestamp 1677592792
<< locali >>
rect 61 1747 69 1781
rect 103 1747 111 1781
rect 61 17 111 1747
rect 577 1747 585 1781
rect 619 1747 627 1781
rect 405 1495 413 1529
rect 447 1495 455 1529
rect 61 -17 69 17
rect 103 -17 111 17
rect 577 17 627 1747
rect 1093 1495 1101 1529
rect 1135 1495 1143 1529
rect 577 -17 585 17
rect 619 -17 627 17
<< viali >>
rect 69 1747 103 1781
rect 585 1747 619 1781
rect 413 1495 447 1529
rect 69 -17 103 17
rect 1101 1495 1135 1529
rect 585 -17 619 17
<< metal1 >>
rect 52 1790 204 1792
rect 52 1781 146 1790
rect 52 1747 69 1781
rect 103 1747 146 1781
rect 52 1738 146 1747
rect 198 1738 204 1790
rect 52 1736 204 1738
rect 568 1790 720 1792
rect 568 1781 662 1790
rect 568 1747 585 1781
rect 619 1747 662 1781
rect 568 1738 662 1747
rect 714 1738 720 1790
rect 568 1736 720 1738
rect 1172 1790 1408 1792
rect 1172 1738 1178 1790
rect 1230 1738 1350 1790
rect 1402 1738 1408 1790
rect 1172 1736 1408 1738
rect 396 1538 806 1540
rect 396 1529 748 1538
rect 396 1495 413 1529
rect 447 1495 748 1529
rect 396 1486 748 1495
rect 800 1486 806 1538
rect 396 1484 806 1486
rect 914 1538 1152 1540
rect 914 1486 920 1538
rect 972 1529 1152 1538
rect 972 1495 1101 1529
rect 1135 1495 1152 1529
rect 972 1486 1152 1495
rect 914 1484 1152 1486
rect 54 1286 204 1288
rect 54 1234 60 1286
rect 112 1234 146 1286
rect 198 1234 204 1286
rect 54 1232 204 1234
rect 570 1286 720 1288
rect 570 1234 576 1286
rect 628 1234 662 1286
rect 714 1234 720 1286
rect 570 1232 720 1234
rect 1258 1286 1408 1288
rect 1258 1234 1264 1286
rect 1316 1234 1350 1286
rect 1402 1234 1408 1286
rect 1258 1232 1408 1234
rect 52 26 120 28
rect 52 -26 60 26
rect 112 -26 120 26
rect 52 -28 120 -26
rect 412 -372 466 610
rect 892 560 1002 616
rect 568 26 636 28
rect 568 -26 576 26
rect 628 -26 636 26
rect 568 -28 636 -26
rect 932 -174 1002 560
rect 1088 472 1150 616
rect 2484 474 2582 482
rect 2484 472 2770 474
rect 1088 404 2492 472
rect 2484 402 2492 404
rect 2572 402 2770 472
rect 2484 400 2770 402
rect 2484 386 2582 400
rect 2368 -174 2484 -152
rect 932 -180 2484 -174
rect 932 -260 2380 -180
rect 2368 -262 2380 -260
rect 2466 -262 2484 -180
rect 2368 -288 2484 -262
rect 412 -422 1006 -372
rect 412 -434 1012 -422
rect 412 -438 930 -434
rect 916 -492 930 -438
rect 1000 -492 1012 -434
rect 916 -502 1012 -492
rect 2386 -490 2468 -288
rect 928 -738 998 -502
rect 2386 -560 3292 -490
rect 3202 -684 3292 -560
<< via1 >>
rect 146 1738 198 1790
rect 662 1738 714 1790
rect 1178 1738 1230 1790
rect 1350 1738 1402 1790
rect 748 1486 800 1538
rect 920 1486 972 1538
rect 60 1234 112 1286
rect 146 1234 198 1286
rect 576 1234 628 1286
rect 662 1234 714 1286
rect 1264 1234 1316 1286
rect 1350 1234 1402 1286
rect 60 17 112 26
rect 60 -17 69 17
rect 69 -17 103 17
rect 103 -17 112 17
rect 60 -26 112 -17
rect 576 17 628 26
rect 576 -17 585 17
rect 585 -17 619 17
rect 619 -17 628 17
rect 576 -26 628 -17
rect 2492 402 2572 472
rect 2380 -262 2466 -180
rect 930 -492 1000 -434
<< metal2 >>
rect 58 1792 114 1801
rect 58 1286 114 1736
rect 144 1790 200 1796
rect 144 1738 146 1790
rect 198 1738 200 1790
rect 144 1732 200 1738
rect 574 1792 630 1801
rect 230 1540 286 1549
rect 230 1475 286 1484
rect 58 1234 60 1286
rect 112 1234 114 1286
rect 58 1228 114 1234
rect 144 1286 200 1292
rect 144 1234 146 1286
rect 198 1234 200 1286
rect 144 1228 200 1234
rect 574 1286 630 1736
rect 660 1790 716 1796
rect 660 1738 662 1790
rect 714 1738 716 1790
rect 660 1732 716 1738
rect 1176 1790 1232 1796
rect 1176 1738 1178 1790
rect 1230 1738 1232 1790
rect 746 1538 802 1544
rect 746 1486 748 1538
rect 800 1486 802 1538
rect 746 1480 802 1486
rect 918 1540 974 1549
rect 918 1475 974 1484
rect 574 1234 576 1286
rect 628 1234 630 1286
rect 574 1228 630 1234
rect 660 1286 716 1292
rect 660 1234 662 1286
rect 714 1234 716 1286
rect 660 1228 716 1234
rect 58 28 114 48
rect 58 -37 114 -28
rect 574 28 630 48
rect 574 -37 630 -28
rect 1176 28 1232 1738
rect 1262 1792 1318 1801
rect 1262 1286 1318 1736
rect 1348 1790 1404 1796
rect 1348 1738 1350 1790
rect 1402 1738 1404 1790
rect 1348 1732 1404 1738
rect 1262 1234 1264 1286
rect 1316 1234 1318 1286
rect 1262 1228 1318 1234
rect 1348 1286 1404 1292
rect 1348 1234 1350 1286
rect 1402 1234 1404 1286
rect 1348 1228 1404 1234
rect 2484 474 2582 482
rect 2484 472 2770 474
rect 2484 402 2492 472
rect 2572 468 2770 472
rect 2572 408 2700 468
rect 2758 408 2770 468
rect 2572 402 2770 408
rect 2484 400 2770 402
rect 2484 386 2582 400
rect 1176 -37 1232 -28
rect 2368 -180 2484 -152
rect 2368 -262 2380 -180
rect 2466 -262 2484 -180
rect 2368 -288 2484 -262
rect 916 -434 1012 -422
rect 916 -492 930 -434
rect 1000 -492 1012 -434
rect 916 -502 1012 -492
rect 2386 -490 2468 -288
rect 928 -670 998 -502
rect 2386 -560 3292 -490
rect 928 -726 938 -670
rect 994 -726 998 -670
rect 3202 -608 3292 -560
rect 3202 -674 3218 -608
rect 3274 -674 3292 -608
rect 3202 -684 3292 -674
rect 928 -738 998 -726
<< via2 >>
rect 58 1736 114 1792
rect 574 1736 630 1792
rect 230 1484 286 1540
rect 918 1538 974 1540
rect 918 1486 920 1538
rect 920 1486 972 1538
rect 972 1486 974 1538
rect 918 1484 974 1486
rect 58 26 114 28
rect 58 -26 60 26
rect 60 -26 112 26
rect 112 -26 114 26
rect 58 -28 114 -26
rect 574 26 630 28
rect 574 -26 576 26
rect 576 -26 628 26
rect 628 -26 630 26
rect 574 -28 630 -26
rect 1262 1736 1318 1792
rect 2700 408 2758 468
rect 1176 -28 1232 28
rect 938 -726 994 -670
rect 3218 -674 3274 -608
<< metal3 >>
rect -80 1796 1842 1844
rect -80 1792 1730 1796
rect -80 1736 58 1792
rect 114 1736 574 1792
rect 630 1736 1262 1792
rect 1318 1736 1730 1792
rect -80 1732 1730 1736
rect 1794 1732 1842 1796
rect -80 1684 1842 1732
rect 225 1540 979 1592
rect 225 1484 230 1540
rect 286 1484 918 1540
rect 974 1484 979 1540
rect 225 1432 979 1484
rect 2748 514 8644 5402
rect 2668 468 8644 514
rect 2668 408 2700 468
rect 2758 408 8644 468
rect 2668 340 8644 408
rect -80 64 1842 80
rect -80 -42 -70 64
rect 36 28 1842 64
rect 36 -28 58 28
rect 114 -28 574 28
rect 630 -28 1176 28
rect 1232 -28 1842 28
rect 36 -42 1842 -28
rect -80 -80 1842 -42
rect 2748 -388 8644 340
rect 3168 -608 3322 -582
rect 3168 -634 3218 -608
rect -3198 -670 2698 -644
rect -3198 -726 938 -670
rect 994 -726 2698 -670
rect -3198 -6434 2698 -726
rect 2836 -674 3218 -634
rect 3274 -634 3322 -608
rect 3274 -674 8732 -634
rect 2836 -6424 8732 -674
<< via3 >>
rect 1730 1732 1794 1796
rect -70 -42 36 64
<< mimcap >>
rect 2798 1092 8592 5338
rect 2798 286 3388 1092
rect 4452 286 8592 1092
rect 2798 -310 8592 286
rect -3146 -972 2648 -748
rect -3146 -1778 1290 -972
rect 2354 -1778 2648 -972
rect -3146 -6396 2648 -1778
rect 2898 -1034 8692 -720
rect 2898 -1840 3186 -1034
rect 4250 -1840 8692 -1034
rect 2898 -6368 8692 -1840
<< mimcapcontact >>
rect 3388 286 4452 1092
rect 1290 -1778 2354 -972
rect 3186 -1840 4250 -1034
<< metal4 >>
rect -118 64 118 3024
rect -118 -42 -70 64
rect 36 -42 118 64
rect -118 -1258 118 -42
rect 1644 1796 1880 1882
rect 1644 1732 1730 1796
rect 1794 1732 1880 1796
rect 1644 -118 1880 1732
rect 3356 1092 4472 1104
rect 3356 286 3388 1092
rect 4452 286 4472 1092
rect 3356 258 4472 286
rect 1270 -972 2386 -956
rect 1270 -1258 1290 -972
rect -118 -1442 1290 -1258
rect 1270 -1778 1290 -1442
rect 2354 -1276 2386 -972
rect 3640 -1016 3914 258
rect 3164 -1034 4280 -1016
rect 3164 -1276 3186 -1034
rect 2354 -1460 3186 -1276
rect 2354 -1778 2386 -1460
rect 1270 -1802 2386 -1778
rect 3164 -1840 3186 -1460
rect 4250 -1840 4280 -1034
rect 3164 -1862 4280 -1840
use INV_21850877_PG0_0_0_1677466712  INV_21850877_PG0_0_0_1677466712_0
timestamp 1677466831
transform -1 0 516 0 1 0
box 0 30 516 3024
use STAGE2_INV_27873531_PG0_0_0_1677466713  STAGE2_INV_27873531_PG0_0_0_1677466713_0
timestamp 1677466831
transform -1 0 1548 0 1 0
box 0 30 1032 3024
<< labels >>
rlabel metal4 -76 836 -76 836 1 VN
port 1 n
rlabel metal4 1758 642 1758 642 1 VP
port 2 n
rlabel metal1 948 526 948 526 1 Y
port 3 n
<< end >>
