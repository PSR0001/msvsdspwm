magic
tech sky130A
magscale 1 2
timestamp 1678383033
<< locali >>
rect 61 1579 69 1613
rect 103 1579 111 1613
rect 61 1445 111 1579
rect 61 1411 69 1445
rect 103 1411 111 1445
<< viali >>
rect 69 1579 103 1613
rect 69 1411 103 1445
<< metal1 >>
rect 226 2462 290 2464
rect 226 2410 232 2462
rect 284 2410 290 2462
rect 226 2408 290 2410
rect 52 1613 120 1624
rect 52 1579 69 1613
rect 103 1579 120 1613
rect 52 1568 120 1579
rect 52 1445 120 1456
rect 52 1411 69 1445
rect 103 1411 120 1445
rect 52 1400 120 1411
rect 226 614 290 616
rect 226 562 232 614
rect 284 562 290 614
rect 226 560 290 562
<< via1 >>
rect 232 2410 284 2462
rect 232 562 284 614
<< metal2 >>
rect 230 2462 286 2468
rect 230 2410 232 2462
rect 284 2410 286 2462
rect 230 614 286 2410
rect 230 562 232 614
rect 284 562 286 614
rect 230 556 286 562
use NMOS_S_94657632_X1_Y1_1678382966_1678382967  NMOS_S_94657632_X1_Y1_1678382966_1678382967_0
timestamp 1678383033
transform 1 0 0 0 -1 1512
box 52 56 395 1482
use PMOS_S_13339638_X1_Y1_1678382967_1678382967  PMOS_S_13339638_X1_Y1_1678382967_1678382967_0
timestamp 1678383033
transform 1 0 0 0 1 1512
box 0 0 516 1512
<< end >>
