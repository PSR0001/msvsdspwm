module ANALOG( input VN, input VY, output reg Y);  
  
@@ @np dummy verilog code


endmodule