magic
tech sky130A
magscale 1 2
timestamp 1677523798
<< error_p >>
rect 19 165 77 171
rect 19 131 31 165
rect 19 125 77 131
rect -77 -131 -19 -125
rect -77 -165 -65 -131
rect -77 -171 -19 -165
<< nwell >>
rect -263 -303 263 303
<< pmos >>
rect -63 -84 -33 84
rect 33 -84 63 84
<< pdiff >>
rect -125 72 -63 84
rect -125 -72 -113 72
rect -79 -72 -63 72
rect -125 -84 -63 -72
rect -33 72 33 84
rect -33 -72 -17 72
rect 17 -72 33 72
rect -33 -84 33 -72
rect 63 72 125 84
rect 63 -72 79 72
rect 113 -72 125 72
rect 63 -84 125 -72
<< pdiffc >>
rect -113 -72 -79 72
rect -17 -72 17 72
rect 79 -72 113 72
<< nsubdiff >>
rect -227 233 -131 267
rect 131 233 227 267
rect -227 171 -193 233
rect 193 171 227 233
rect -227 -233 -193 -171
rect 193 -233 227 -171
rect -227 -267 -131 -233
rect 131 -267 227 -233
<< nsubdiffcont >>
rect -131 233 131 267
rect -227 -171 -193 171
rect 193 -171 227 171
rect -131 -267 131 -233
<< poly >>
rect 15 165 81 181
rect 15 131 31 165
rect 65 131 81 165
rect 15 115 81 131
rect -63 84 -33 110
rect 33 84 63 115
rect -63 -115 -33 -84
rect 33 -110 63 -84
rect -81 -131 -15 -115
rect -81 -165 -65 -131
rect -31 -165 -15 -131
rect -81 -181 -15 -165
<< polycont >>
rect 31 131 65 165
rect -65 -165 -31 -131
<< locali >>
rect -227 233 -131 267
rect 131 233 227 267
rect -227 171 -193 233
rect 193 171 227 233
rect 15 131 31 165
rect 65 131 81 165
rect -113 72 -79 88
rect -113 -88 -79 -72
rect -17 72 17 88
rect -17 -88 17 -72
rect 79 72 113 88
rect 79 -88 113 -72
rect -81 -165 -65 -131
rect -31 -165 -15 -131
rect -227 -233 -193 -171
rect 193 -233 227 -171
rect -227 -267 -131 -233
rect 131 -267 227 -233
<< viali >>
rect 31 131 65 165
rect -113 -72 -79 72
rect -17 -72 17 72
rect 79 -72 113 72
rect -65 -165 -31 -131
<< metal1 >>
rect 19 165 77 171
rect 19 131 31 165
rect 65 131 77 165
rect 19 125 77 131
rect -119 72 -73 84
rect -119 -72 -113 72
rect -79 -72 -73 72
rect -119 -84 -73 -72
rect -23 72 23 84
rect -23 -72 -17 72
rect 17 -72 23 72
rect -23 -84 23 -72
rect 73 72 119 84
rect 73 -72 79 72
rect 113 -72 119 72
rect 73 -84 119 -72
rect -77 -131 -19 -125
rect -77 -165 -65 -131
rect -31 -165 -19 -131
rect -77 -171 -19 -165
<< properties >>
string FIXED_BBOX -210 -250 210 250
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 0.84 l 0.15 m 1 nf 2 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
