* NGSPICE file created from Function_Sky130.ext - technology: sky130A

.subckt sky130_fd_pr__pfet_01v8_XGS3BL a_n73_n100# a_15_n100# w_n211_n319# a_n33_n197#
+ VSUBS
X0 a_15_n100# a_n33_n197# a_n73_n100# w_n211_n319# sky130_fd_pr__pfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
C0 a_n73_n100# a_n33_n197# 0.03fF
C1 a_n73_n100# a_15_n100# 0.16fF
C2 a_n33_n197# a_15_n100# 0.03fF
C3 a_n73_n100# w_n211_n319# 0.09fF
C4 w_n211_n319# a_n33_n197# 0.26fF
C5 w_n211_n319# a_15_n100# 0.06fF
C6 a_15_n100# VSUBS 0.02fF
C7 a_n73_n100# VSUBS 0.02fF
C8 a_n33_n197# VSUBS 0.05fF
C9 w_n211_n319# VSUBS 1.07fF
.ends

.subckt sky130_fd_pr__nfet_01v8_648S5X a_n73_n100# a_n33_n188# a_15_n100# a_n175_n274#
X0 a_15_n100# a_n33_n188# a_n73_n100# a_n175_n274# sky130_fd_pr__nfet_01v8 ad=2.9e+11p pd=2.58e+06u as=2.9e+11p ps=2.58e+06u w=1e+06u l=150000u
C0 a_15_n100# a_n73_n100# 0.16fF
C1 a_15_n100# a_n33_n188# 0.03fF
C2 a_n33_n188# a_n73_n100# 0.03fF
C3 a_15_n100# a_n175_n274# 0.08fF
C4 a_n73_n100# a_n175_n274# 0.11fF
C5 a_n33_n188# a_n175_n274# 0.30fF
.ends

.subckt Function_Sky130 A C E F D B Y VDD GND
XXM12 m1_738_2130# m1_2538_2132# w_n208_1792# D VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM1 Y A m1_136_1220# VSUBS sky130_fd_pr__nfet_01v8_648S5X
XXM2 m1_136_1220# C Y VSUBS sky130_fd_pr__nfet_01v8_648S5X
XXM3 Y E m1_1334_1224# VSUBS sky130_fd_pr__nfet_01v8_648S5X
XXM4 m1_1334_1224# F GND VSUBS sky130_fd_pr__nfet_01v8_648S5X
XXM5 m1_136_1220# B GND VSUBS sky130_fd_pr__nfet_01v8_648S5X
XXM6 GND D m1_136_1220# VSUBS sky130_fd_pr__nfet_01v8_648S5X
XXM7 m1_738_2130# Y w_n208_1792# E VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM8 Y m1_738_2130# w_n208_1792# F VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM9 VDD m1_136_2130# w_n208_1792# A VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM10 m1_136_2130# m1_738_2130# w_n208_1792# C VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
XXM11 m1_2538_2132# VDD w_n208_1792# B VSUBS sky130_fd_pr__pfet_01v8_XGS3BL
C0 B m1_1334_1224# 0.00fF
C1 F m1_738_2130# 0.15fF
C2 m1_136_1220# m1_2538_2132# 0.00fF
C3 D m1_2538_2132# 0.10fF
C4 A m1_738_2130# 0.00fF
C5 Y m1_136_1220# 0.29fF
C6 D Y 0.17fF
C7 m1_1334_1224# GND 0.08fF
C8 C GND 0.03fF
C9 B GND 0.16fF
C10 m1_136_2130# C 0.10fF
C11 m1_1334_1224# E 0.10fF
C12 m1_136_1220# w_n208_1792# 0.42fF
C13 E C 0.12fF
C14 D w_n208_1792# 0.35fF
C15 VDD m1_136_1220# 0.00fF
C16 D VDD 0.02fF
C17 F m1_136_1220# 0.07fF
C18 D F 0.12fF
C19 A m1_136_1220# 0.20fF
C20 m1_738_2130# m1_136_1220# 0.01fF
C21 m1_1334_1224# Y 0.08fF
C22 D m1_738_2130# 0.12fF
C23 Y C 0.27fF
C24 B m1_2538_2132# 0.10fF
C25 E GND 0.03fF
C26 B Y 0.15fF
C27 m1_136_2130# E 0.00fF
C28 m1_1334_1224# w_n208_1792# 0.00fF
C29 C w_n208_1792# 0.25fF
C30 Y GND 0.22fF
C31 C VDD 0.02fF
C32 m1_1334_1224# F 0.10fF
C33 B w_n208_1792# 0.24fF
C34 F C 0.00fF
C35 m1_136_2130# Y 0.05fF
C36 E m1_2538_2132# 0.00fF
C37 B VDD 0.13fF
C38 m1_1334_1224# A 0.00fF
C39 D m1_136_1220# 0.27fF
C40 Y E 0.38fF
C41 C A 0.11fF
C42 B F 0.00fF
C43 C m1_738_2130# 0.11fF
C44 B m1_738_2130# 0.00fF
C45 GND w_n208_1792# 0.09fF
C46 GND VDD 0.00fF
C47 Y m1_2538_2132# 0.05fF
C48 m1_136_2130# w_n208_1792# 0.19fF
C49 F GND 0.14fF
C50 m1_136_2130# VDD 0.05fF
C51 E w_n208_1792# 0.31fF
C52 A GND 0.04fF
C53 m1_136_2130# F 0.00fF
C54 E VDD 0.00fF
C55 F E 0.12fF
C56 m1_136_2130# A 0.09fF
C57 m1_136_2130# m1_738_2130# 0.00fF
C58 m1_2538_2132# w_n208_1792# 0.21fF
C59 E A 0.00fF
C60 m1_1334_1224# m1_136_1220# 0.12fF
C61 VDD m1_2538_2132# 0.05fF
C62 m1_1334_1224# D 0.00fF
C63 E m1_738_2130# 0.15fF
C64 C m1_136_1220# 0.23fF
C65 Y w_n208_1792# 4.06fF
C66 Y VDD 0.05fF
C67 F m1_2538_2132# 0.00fF
C68 B m1_136_1220# 0.17fF
C69 B D 0.12fF
C70 Y F 0.28fF
C71 m1_738_2130# m1_2538_2132# 0.00fF
C72 Y A 0.26fF
C73 Y m1_738_2130# 0.18fF
C74 GND m1_136_1220# 4.80fF
C75 D GND 0.14fF
C76 VDD w_n208_1792# 5.57fF
C77 F w_n208_1792# 0.29fF
C78 m1_136_2130# m1_136_1220# 0.00fF
C79 F VDD 0.00fF
C80 E m1_136_1220# 0.06fF
C81 D E 0.00fF
C82 A w_n208_1792# 0.15fF
C83 m1_1334_1224# C 0.00fF
C84 A VDD 0.13fF
C85 m1_738_2130# w_n208_1792# 1.59fF
C86 m1_738_2130# VDD 0.81fF
C87 m1_738_2130# VSUBS -1.43fF
C88 m1_136_2130# VSUBS -0.03fF
C89 VDD VSUBS -5.27fF
C90 w_n208_1792# VSUBS 10.28fF
C91 D VSUBS 0.09fF
C92 B VSUBS 0.43fF
C93 GND VSUBS 0.18fF
C94 F VSUBS 0.19fF
C95 m1_1334_1224# VSUBS 0.27fF
C96 E VSUBS 0.16fF
C97 C VSUBS 0.22fF
C98 m1_136_1220# VSUBS -1.33fF
C99 Y VSUBS -6.17fF
C100 A VSUBS 0.47fF
C101 m1_2538_2132# VSUBS -0.25fF
.ends



Vdd VDD GND 1.8
.save i(vdd)
Vdd1 A GND pulse(0 1.8 0.1n 10p 10p 1n 2n)
.save i(vdd1)
Vdd2 B GND pulse(0 1.8 0.2n 10p 10p 1n 2n)
.save i(vdd2)
Vdd3 C GND pulse(0 1.8 0.3n 10p 10p 1n 2n)
.save i(vdd3)
Vdd4 D GND pulse(0 1.8 0.4n 10p 10p 1n 2n)
.save i(vdd4)
Vdd5 E GND pulse(0 1.8 0.5n 10p 10p 1n 2n)
.save i(vdd5)
Vdd6 F GND pulse(0 1.8 0.6n 10p 10p 1n 2n)
.save i(vdd6)
X1 F E D C B A  Y VDD GND  Function_Sky130
**** begin user architecture code


.lib ~/open_pdks/sources/sky130-pdk/libraries/sky130_fd_pr/latest/models/sky130.lib.spice tt
.control
save all
tran 10p 4n
plot y
.endc
