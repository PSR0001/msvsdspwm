magic
tech sky130A
magscale 1 2
timestamp 1677862335
<< metal1 >>
rect 312 2462 376 2464
rect 312 2410 318 2462
rect 370 2410 376 2462
rect 312 2408 376 2410
rect 226 1622 290 1624
rect 226 1570 232 1622
rect 284 1570 290 1622
rect 226 1568 290 1570
rect 226 1454 290 1456
rect 226 1402 232 1454
rect 284 1402 290 1454
rect 226 1400 290 1402
rect 312 614 376 616
rect 312 562 318 614
rect 370 562 376 614
rect 312 560 376 562
<< via1 >>
rect 318 2410 370 2462
rect 232 1570 284 1622
rect 232 1402 284 1454
rect 318 562 370 614
<< metal2 >>
rect 316 2462 372 2468
rect 316 2410 318 2462
rect 370 2410 372 2462
rect 230 1622 286 1628
rect 230 1570 232 1622
rect 284 1570 286 1622
rect 230 1454 286 1570
rect 230 1402 232 1454
rect 284 1402 286 1454
rect 230 1396 286 1402
rect 316 614 372 2410
rect 316 562 318 614
rect 370 562 372 614
rect 316 556 372 562
use NMOS_S_4459928_X5_Y1_1677862245_1677862246  NMOS_S_4459928_X5_Y1_1677862245_1677862246_0
timestamp 1677862335
transform 1 0 0 0 -1 1512
box 121 56 1083 1482
use PMOS_S_62253992_X5_Y1_1677862246_1677862246  PMOS_S_62253992_X5_Y1_1677862246_1677862246_0
timestamp 1677862335
transform 1 0 0 0 1 1512
box 0 0 1204 1512
<< end >>
