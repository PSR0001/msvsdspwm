magic
tech sky130A
magscale 1 2
timestamp 1677519681
<< locali >>
rect 61 1579 69 1613
rect 103 1579 111 1613
rect 61 1445 111 1579
rect 61 1411 69 1445
rect 103 1411 111 1445
<< viali >>
rect 69 1579 103 1613
rect 69 1411 103 1445
<< metal1 >>
rect 54 2462 118 2464
rect 54 2410 60 2462
rect 112 2410 118 2462
rect 54 2408 118 2410
rect 52 1613 120 1624
rect 52 1579 69 1613
rect 103 1579 120 1613
rect 52 1568 120 1579
rect 52 1445 120 1456
rect 52 1411 69 1445
rect 103 1411 120 1445
rect 52 1400 120 1411
rect 54 614 118 616
rect 54 562 60 614
rect 112 562 118 614
rect 54 560 118 562
<< via1 >>
rect 60 2410 112 2462
rect 60 562 112 614
<< metal2 >>
rect 58 2462 114 2468
rect 58 2410 60 2462
rect 112 2410 114 2462
rect 58 614 114 2410
rect 58 562 60 614
rect 112 562 114 614
rect 58 556 114 562
use NMOS_S_25628869_X1_Y1_1677518941_1677518943  NMOS_S_25628869_X1_Y1_1677518941_1677518943_0
timestamp 1677519681
transform 1 0 0 0 -1 1512
box 52 56 395 1482
use PMOS_S_89421238_X1_Y1_1677518942_1677518943  PMOS_S_89421238_X1_Y1_1677518942_1677518943_0
timestamp 1677519681
transform 1 0 0 0 1 1512
box 0 0 516 1512
<< end >>
