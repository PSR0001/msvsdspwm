magic
tech sky130A
magscale 1 2
timestamp 1677466831
<< nwell >>
rect 0 0 516 1512
<< pmos >>
rect 200 399 230 735
rect 286 399 316 735
<< pdiff >>
rect 147 585 200 735
rect 147 551 155 585
rect 189 551 200 585
rect 147 517 200 551
rect 147 483 155 517
rect 189 483 200 517
rect 147 449 200 483
rect 147 415 155 449
rect 189 415 200 449
rect 147 399 200 415
rect 230 585 286 735
rect 230 551 241 585
rect 275 551 286 585
rect 230 517 286 551
rect 230 483 241 517
rect 275 483 286 517
rect 230 449 286 483
rect 230 415 241 449
rect 275 415 286 449
rect 230 399 286 415
rect 316 585 369 735
rect 316 551 327 585
rect 361 551 369 585
rect 316 517 369 551
rect 316 483 327 517
rect 361 483 369 517
rect 316 449 369 483
rect 316 415 327 449
rect 361 415 369 449
rect 316 399 369 415
<< pdiffc >>
rect 155 551 189 585
rect 155 483 189 517
rect 155 415 189 449
rect 241 551 275 585
rect 241 483 275 517
rect 241 415 275 449
rect 327 551 361 585
rect 327 483 361 517
rect 327 415 361 449
<< nsubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
<< nsubdiffcont >>
rect 241 1327 275 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 735 230 897
rect 286 735 316 897
rect 200 252 230 399
rect 286 252 316 399
<< polycont >>
rect 241 907 275 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 147 585 197 773
rect 147 551 155 585
rect 189 551 197 585
rect 147 517 197 551
rect 147 483 155 517
rect 189 483 197 517
rect 147 449 197 483
rect 147 415 155 449
rect 189 415 197 449
rect 147 185 197 415
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 585 283 773
rect 233 551 241 585
rect 275 551 283 585
rect 233 517 283 551
rect 233 483 241 517
rect 275 483 283 517
rect 233 449 283 483
rect 233 415 241 449
rect 275 415 283 449
rect 233 101 283 415
rect 233 67 241 101
rect 275 67 283 101
rect 319 585 369 773
rect 319 551 327 585
rect 361 551 369 585
rect 319 517 369 551
rect 319 483 327 517
rect 361 483 369 517
rect 319 449 369 483
rect 319 415 327 449
rect 361 415 369 449
rect 319 185 369 415
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
<< viali >>
rect 241 1327 275 1361
rect 241 907 275 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
<< metal1 >>
rect 138 1370 378 1372
rect 138 1361 318 1370
rect 138 1327 241 1361
rect 275 1327 318 1361
rect 138 1318 318 1327
rect 370 1318 378 1370
rect 138 1316 378 1318
rect 52 941 292 952
rect 52 907 241 941
rect 275 907 292 941
rect 52 896 292 907
rect 138 194 378 196
rect 138 185 318 194
rect 138 151 155 185
rect 189 151 318 185
rect 138 142 318 151
rect 370 142 378 194
rect 138 140 378 142
rect 52 101 292 112
rect 52 67 241 101
rect 275 67 292 101
rect 52 56 292 67
<< via1 >>
rect 318 1318 370 1370
rect 318 185 370 194
rect 318 151 327 185
rect 327 151 361 185
rect 361 151 370 185
rect 318 142 370 151
<< metal2 >>
rect 316 1370 372 1376
rect 316 1318 318 1370
rect 370 1318 372 1370
rect 316 194 372 1318
rect 316 142 318 194
rect 370 142 372 194
rect 316 136 372 142
<< end >>
