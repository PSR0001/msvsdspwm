magic
tech sky130A
magscale 1 2
timestamp 1676459712
<< locali >>
rect 921 1579 929 1613
rect 963 1579 971 1613
rect 921 1445 971 1579
rect 921 1411 929 1445
rect 963 1411 971 1445
rect 1093 1495 1101 1529
rect 1135 1495 1143 1529
rect 1093 1445 1143 1495
rect 1093 1411 1101 1445
rect 1135 1411 1143 1445
rect 2813 571 2821 605
rect 2855 571 2863 605
rect 2813 521 2863 571
rect 2813 487 2821 521
rect 2855 487 2863 521
<< viali >>
rect 929 1579 963 1613
rect 929 1411 963 1445
rect 1101 1495 1135 1529
rect 1101 1411 1135 1445
rect 2821 571 2855 605
rect 2821 487 2855 521
<< metal1 >>
rect 1806 2408 1978 2464
rect 2838 2408 3010 2464
rect 912 1613 1634 1624
rect 912 1579 929 1613
rect 963 1579 1634 1613
rect 912 1568 1634 1579
rect 1774 1622 1838 1624
rect 1774 1570 1780 1622
rect 1832 1570 1838 1622
rect 1774 1568 1838 1570
rect 1946 1622 2010 1624
rect 1946 1570 1952 1622
rect 2004 1570 2010 1622
rect 1946 1568 2010 1570
rect 2150 1568 2666 1624
rect 2978 1622 3042 1624
rect 2978 1570 2984 1622
rect 3036 1570 3042 1622
rect 2978 1568 3042 1570
rect 312 1538 1152 1540
rect 312 1486 318 1538
rect 370 1529 1152 1538
rect 370 1495 1101 1529
rect 1135 1495 1152 1529
rect 370 1486 1152 1495
rect 312 1484 1152 1486
rect 1516 1538 1752 1540
rect 1516 1486 1522 1538
rect 1574 1486 1694 1538
rect 1746 1486 1752 1538
rect 1516 1484 1752 1486
rect 2462 1538 2612 1540
rect 2462 1486 2468 1538
rect 2520 1486 2554 1538
rect 2606 1486 2612 1538
rect 2462 1484 2612 1486
rect 3064 1538 3300 1540
rect 3064 1486 3070 1538
rect 3122 1486 3242 1538
rect 3294 1486 3300 1538
rect 3064 1484 3300 1486
rect 258 1400 774 1456
rect 912 1445 980 1456
rect 912 1411 929 1445
rect 963 1411 980 1445
rect 912 1400 980 1411
rect 1084 1445 1152 1456
rect 1084 1411 1101 1445
rect 1135 1411 1152 1445
rect 1084 1400 1152 1411
rect 1774 1454 1838 1456
rect 1774 1402 1780 1454
rect 1832 1402 1838 1454
rect 1774 1400 1838 1402
rect 2204 1454 2268 1456
rect 2204 1402 2210 1454
rect 2262 1402 2268 1454
rect 2204 1400 2268 1402
rect 2634 1454 2838 1456
rect 2634 1402 2640 1454
rect 2692 1402 2838 1454
rect 2634 1400 2838 1402
rect 2978 1454 3042 1456
rect 2978 1402 2984 1454
rect 3036 1402 3042 1454
rect 2978 1400 3042 1402
rect 2462 1370 2526 1372
rect 2462 1318 2468 1370
rect 2520 1318 2526 1370
rect 2462 1316 2526 1318
rect 946 560 1118 616
rect 1978 560 2150 616
rect 2804 605 2872 616
rect 2804 571 2821 605
rect 2855 571 2872 605
rect 2804 560 2872 571
rect 2494 521 2872 532
rect 2494 487 2821 521
rect 2855 487 2872 521
rect 2494 476 2872 487
rect 312 278 720 280
rect 312 226 318 278
rect 370 226 662 278
rect 714 226 720 278
rect 312 224 720 226
rect 1344 278 3128 280
rect 1344 226 1350 278
rect 1402 226 3070 278
rect 3122 226 3128 278
rect 1344 224 3128 226
<< via1 >>
rect 1780 1570 1832 1622
rect 1952 1570 2004 1622
rect 2984 1570 3036 1622
rect 318 1486 370 1538
rect 1522 1486 1574 1538
rect 1694 1486 1746 1538
rect 2468 1486 2520 1538
rect 2554 1486 2606 1538
rect 3070 1486 3122 1538
rect 3242 1486 3294 1538
rect 1780 1402 1832 1454
rect 2210 1402 2262 1454
rect 2640 1402 2692 1454
rect 2984 1402 3036 1454
rect 2468 1318 2520 1370
rect 318 226 370 278
rect 662 226 714 278
rect 1350 226 1402 278
rect 3070 226 3122 278
<< metal2 >>
rect 316 1538 372 1568
rect 316 1486 318 1538
rect 370 1486 372 1538
rect 316 1480 372 1486
rect 660 1540 716 1549
rect 660 1344 716 1484
rect 1520 1538 1576 1680
rect 1778 1622 1834 1628
rect 1778 1570 1780 1622
rect 1832 1570 1834 1622
rect 1520 1486 1522 1538
rect 1574 1486 1576 1538
rect 1520 1480 1576 1486
rect 1692 1538 1748 1544
rect 1692 1486 1694 1538
rect 1746 1486 1748 1538
rect 1692 1344 1748 1486
rect 1778 1454 1834 1570
rect 1950 1622 2006 1628
rect 1950 1570 1952 1622
rect 2004 1570 2006 1622
rect 1950 1540 2006 1570
rect 1950 1475 2006 1484
rect 1778 1402 1780 1454
rect 1832 1402 1834 1454
rect 1778 1396 1834 1402
rect 2208 1454 2264 1680
rect 2208 1402 2210 1454
rect 2262 1402 2264 1454
rect 2208 1396 2264 1402
rect 2466 1538 2522 1544
rect 2466 1486 2468 1538
rect 2520 1486 2522 1538
rect 2466 1370 2522 1486
rect 2552 1538 2608 1680
rect 2552 1486 2554 1538
rect 2606 1486 2608 1538
rect 2552 1480 2608 1486
rect 2982 1622 3038 1628
rect 2982 1570 2984 1622
rect 3036 1570 3038 1622
rect 2466 1318 2468 1370
rect 2520 1318 2522 1370
rect 2466 1312 2522 1318
rect 2638 1454 2694 1460
rect 2638 1402 2640 1454
rect 2692 1402 2694 1454
rect 1692 1288 1748 1297
rect 1692 1223 1748 1232
rect 2638 1288 2694 1402
rect 2982 1454 3038 1570
rect 2982 1402 2984 1454
rect 3036 1402 3038 1454
rect 2982 1396 3038 1402
rect 3068 1538 3124 1544
rect 3068 1486 3070 1538
rect 3122 1486 3124 1538
rect 3068 1344 3124 1486
rect 3240 1538 3296 1680
rect 3240 1486 3242 1538
rect 3294 1486 3296 1538
rect 3240 1480 3296 1486
rect 2638 1223 2694 1232
rect 316 278 372 284
rect 316 226 318 278
rect 370 226 372 278
rect 316 220 372 226
rect 660 278 716 284
rect 660 226 662 278
rect 714 226 716 278
rect 660 220 716 226
rect 1348 278 1404 284
rect 1348 226 1350 278
rect 1402 226 1404 278
rect 1348 220 1404 226
rect 3068 278 3124 284
rect 3068 226 3070 278
rect 3122 226 3124 278
rect 3068 220 3124 226
<< via2 >>
rect 660 1484 716 1540
rect 1950 1484 2006 1540
rect 1692 1232 1748 1288
rect 2638 1232 2694 1288
<< metal3 >>
rect 655 1540 2011 1592
rect 655 1484 660 1540
rect 716 1484 1950 1540
rect 2006 1484 2011 1540
rect 655 1432 2011 1484
rect 1687 1288 2699 1340
rect 1687 1232 1692 1288
rect 1748 1232 2638 1288
rect 2694 1232 2699 1288
rect 1687 1180 2699 1232
use DP_PMOS_90543401_X1_Y1_1676446839  DP_PMOS_90543401_X1_Y1_1676446839_0
timestamp 1676458286
transform 1 0 2064 0 -1 1512
box 0 0 688 1512
use INV_6743645_0_0_1676446838  INV_6743645_0_0_1676446838_0
timestamp 1676458286
transform -1 0 516 0 -1 3024
box 0 30 516 3024
use NMOS_S_96839798_X1_Y1_1676446840  NMOS_S_96839798_X1_Y1_1676446840_0
timestamp 1676458286
transform -1 0 1892 0 1 1512
box 52 56 395 1482
use NMOS_S_96839798_X1_Y1_1676446840  NMOS_S_96839798_X1_Y1_1676446840_1
timestamp 1676458286
transform -1 0 2064 0 -1 1512
box 52 56 395 1482
use NMOS_S_96839798_X1_Y1_1676446840  NMOS_S_96839798_X1_Y1_1676446840_2
timestamp 1676458286
transform 1 0 1032 0 -1 1512
box 52 56 395 1482
use NMOS_S_96839798_X1_Y1_1676446840  NMOS_S_96839798_X1_Y1_1676446840_3
timestamp 1676458286
transform 1 0 2924 0 1 1512
box 52 56 395 1482
use NMOS_S_96839798_X1_Y1_1676446840  NMOS_S_96839798_X1_Y1_1676446840_4
timestamp 1676458286
transform 1 0 2752 0 -1 1512
box 52 56 395 1482
use PMOS_S_36030836_X1_Y1_1676446841  PMOS_S_36030836_X1_Y1_1676446841_0
timestamp 1676458286
transform -1 0 2924 0 1 1512
box 0 0 516 1512
use PMOS_S_36030836_X1_Y1_1676446841  PMOS_S_36030836_X1_Y1_1676446841_1
timestamp 1676458286
transform 1 0 1892 0 1 1512
box 0 0 516 1512
use PMOS_S_36030836_X1_Y1_1676446841  PMOS_S_36030836_X1_Y1_1676446841_2
timestamp 1676458286
transform -1 0 1032 0 -1 1512
box 0 0 516 1512
<< labels >>
flabel metal1 s 172 588 172 588 0 FreeSerif 0 0 0 0 E
flabel metal1 s 172 1428 172 1428 0 FreeSerif 0 0 0 0 Y
flabel metal1 s 1892 588 1892 588 0 FreeSerif 0 0 0 0 A
flabel metal1 s 2408 504 2408 504 0 FreeSerif 0 0 0 0 B
flabel metal2 s 2580 714 2580 714 0 FreeSerif 0 0 0 0 VDD
flabel metal2 s 1376 756 1376 756 0 FreeSerif 0 0 0 0 VSS
flabel metal1 s 2752 2436 2752 2436 0 FreeSerif 0 0 0 0 D
flabel metal1 s 860 588 860 588 0 FreeSerif 0 0 0 0 F
flabel metal1 s 1720 2436 1720 2436 0 FreeSerif 0 0 0 0 C
<< end >>
