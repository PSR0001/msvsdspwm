MACRO TEST
  ORIGIN 0 0 ;
  FOREIGN TEST 0 0 ;
  SIZE 17.2 BY 15.12 ;
  PIN E
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
      LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
      LAYER M2 ;
        RECT 0.27 2.8 0.59 3.08 ;
      LAYER M3 ;
        RECT 0.29 2.94 0.57 12.18 ;
      LAYER M2 ;
        RECT 0.27 12.04 0.59 12.32 ;
    END
  END E
  PIN Y
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
      LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
      LAYER M2 ;
        RECT 0.27 7 0.59 7.28 ;
      LAYER M1 ;
        RECT 0.305 7.14 0.555 7.98 ;
      LAYER M2 ;
        RECT 0.27 7.84 0.59 8.12 ;
      LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
      LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
      LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
      LAYER M2 ;
        RECT 1.29 7 3.87 7.28 ;
      LAYER M2 ;
        RECT 4.57 7 4.89 7.28 ;
      LAYER M1 ;
        RECT 4.605 7.14 4.855 7.98 ;
      LAYER M2 ;
        RECT 4.73 7.84 8.17 8.12 ;
      LAYER M2 ;
        RECT 8.87 7.84 9.19 8.12 ;
      LAYER M3 ;
        RECT 8.89 7.14 9.17 7.98 ;
      LAYER M2 ;
        RECT 8.87 7 9.19 7.28 ;
    END
  END Y
  PIN A
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
      LAYER M2 ;
        RECT 10.58 2.8 11.78 3.08 ;
      LAYER M2 ;
        RECT 9.89 2.8 10.75 3.08 ;
    END
  END A
  PIN B
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 11.44 2.38 12.64 2.66 ;
      LAYER M2 ;
        RECT 14.02 2.8 15.22 3.08 ;
      LAYER M2 ;
        RECT 12.47 2.38 14.19 2.66 ;
      LAYER M1 ;
        RECT 14.065 2.52 14.315 2.94 ;
      LAYER M2 ;
        RECT 14.03 2.8 14.35 3.08 ;
    END
  END B
  PIN VDD
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 12.76 0.68 13.04 6.46 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
      LAYER M3 ;
        RECT 15.34 0.68 15.62 6.88 ;
      LAYER M3 ;
        RECT 16.2 8.24 16.48 14.44 ;
      LAYER M3 ;
        RECT 6.74 1.075 7.02 1.445 ;
      LAYER M2 ;
        RECT 6.88 1.12 15.48 1.4 ;
      LAYER M3 ;
        RECT 15.34 1.075 15.62 1.445 ;
      LAYER M3 ;
        RECT 15.34 6.72 15.62 7.56 ;
      LAYER M2 ;
        RECT 15.48 7.42 16.34 7.7 ;
      LAYER M3 ;
        RECT 16.2 7.56 16.48 8.4 ;
    END
  END VSS
  PIN D
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 13.16 12.04 14.36 12.32 ;
      LAYER M2 ;
        RECT 14.88 12.04 16.08 12.32 ;
      LAYER M2 ;
        RECT 14.19 12.04 15.05 12.32 ;
    END
  END D
  PIN F
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
      LAYER M2 ;
        RECT 5.42 2.8 6.62 3.08 ;
      LAYER M2 ;
        RECT 4.73 2.8 5.59 3.08 ;
    END
  END F
  PIN C
    DIRECTION INOUT ;
    USE SIGNAL ;
    PORT 
      LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
      LAYER M2 ;
        RECT 9.72 12.04 10.92 12.32 ;
      LAYER M2 ;
        RECT 9.03 12.04 9.89 12.32 ;
    END
  END C
  OBS 
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M2 ;
        RECT 5.42 7 6.62 7.28 ;
  LAYER M3 ;
        RECT 1.58 7.56 1.86 8.4 ;
  LAYER M2 ;
        RECT 1.72 7.42 5.59 7.7 ;
  LAYER M1 ;
        RECT 5.465 7.14 5.715 7.56 ;
  LAYER M2 ;
        RECT 5.43 7 5.75 7.28 ;
  LAYER M1 ;
        RECT 5.465 7.055 5.715 7.225 ;
  LAYER M2 ;
        RECT 5.42 7 5.76 7.28 ;
  LAYER M1 ;
        RECT 5.465 7.475 5.715 7.645 ;
  LAYER M2 ;
        RECT 5.42 7.42 5.76 7.7 ;
  LAYER M2 ;
        RECT 1.56 7.42 1.88 7.7 ;
  LAYER M3 ;
        RECT 1.58 7.4 1.86 7.72 ;
  LAYER M1 ;
        RECT 5.465 7.055 5.715 7.225 ;
  LAYER M2 ;
        RECT 5.42 7 5.76 7.28 ;
  LAYER M1 ;
        RECT 5.465 7.475 5.715 7.645 ;
  LAYER M2 ;
        RECT 5.42 7.42 5.76 7.7 ;
  LAYER M2 ;
        RECT 1.56 7.42 1.88 7.7 ;
  LAYER M3 ;
        RECT 1.58 7.4 1.86 7.72 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M2 ;
        RECT 9.72 7.84 10.92 8.12 ;
  LAYER M2 ;
        RECT 13.16 7.84 14.36 8.12 ;
  LAYER M3 ;
        RECT 1.58 1.075 1.86 1.445 ;
  LAYER M2 ;
        RECT 1.72 1.12 3.44 1.4 ;
  LAYER M3 ;
        RECT 3.3 1.075 3.58 1.445 ;
  LAYER M3 ;
        RECT 3.3 6.72 3.58 7.56 ;
  LAYER M4 ;
        RECT 3.44 7.16 9.89 7.96 ;
  LAYER M3 ;
        RECT 9.75 7.56 10.03 7.98 ;
  LAYER M2 ;
        RECT 9.73 7.84 10.05 8.12 ;
  LAYER M2 ;
        RECT 10.75 7.84 13.33 8.12 ;
  LAYER M2 ;
        RECT 1.56 1.12 1.88 1.4 ;
  LAYER M3 ;
        RECT 1.58 1.1 1.86 1.42 ;
  LAYER M2 ;
        RECT 3.28 1.12 3.6 1.4 ;
  LAYER M3 ;
        RECT 3.3 1.1 3.58 1.42 ;
  LAYER M2 ;
        RECT 1.56 1.12 1.88 1.4 ;
  LAYER M3 ;
        RECT 1.58 1.1 1.86 1.42 ;
  LAYER M2 ;
        RECT 3.28 1.12 3.6 1.4 ;
  LAYER M3 ;
        RECT 3.3 1.1 3.58 1.42 ;
  LAYER M2 ;
        RECT 1.56 1.12 1.88 1.4 ;
  LAYER M3 ;
        RECT 1.58 1.1 1.86 1.42 ;
  LAYER M2 ;
        RECT 3.28 1.12 3.6 1.4 ;
  LAYER M3 ;
        RECT 3.3 1.1 3.58 1.42 ;
  LAYER M2 ;
        RECT 9.73 7.84 10.05 8.12 ;
  LAYER M3 ;
        RECT 9.75 7.82 10.03 8.14 ;
  LAYER M3 ;
        RECT 3.3 7.375 3.58 7.745 ;
  LAYER M4 ;
        RECT 3.275 7.16 3.605 7.96 ;
  LAYER M3 ;
        RECT 9.75 7.375 10.03 7.745 ;
  LAYER M4 ;
        RECT 9.725 7.16 10.055 7.96 ;
  LAYER M2 ;
        RECT 1.56 1.12 1.88 1.4 ;
  LAYER M3 ;
        RECT 1.58 1.1 1.86 1.42 ;
  LAYER M2 ;
        RECT 3.28 1.12 3.6 1.4 ;
  LAYER M3 ;
        RECT 3.3 1.1 3.58 1.42 ;
  LAYER M2 ;
        RECT 9.73 7.84 10.05 8.12 ;
  LAYER M3 ;
        RECT 9.75 7.82 10.03 8.14 ;
  LAYER M3 ;
        RECT 3.3 7.375 3.58 7.745 ;
  LAYER M4 ;
        RECT 3.275 7.16 3.605 7.96 ;
  LAYER M3 ;
        RECT 9.75 7.375 10.03 7.745 ;
  LAYER M4 ;
        RECT 9.725 7.16 10.055 7.96 ;
  LAYER M2 ;
        RECT 1.56 1.12 1.88 1.4 ;
  LAYER M3 ;
        RECT 1.58 1.1 1.86 1.42 ;
  LAYER M2 ;
        RECT 3.28 1.12 3.6 1.4 ;
  LAYER M3 ;
        RECT 3.3 1.1 3.58 1.42 ;
  LAYER M2 ;
        RECT 9.73 7.84 10.05 8.12 ;
  LAYER M3 ;
        RECT 9.75 7.82 10.03 8.14 ;
  LAYER M3 ;
        RECT 3.3 7.375 3.58 7.745 ;
  LAYER M4 ;
        RECT 3.275 7.16 3.605 7.96 ;
  LAYER M3 ;
        RECT 9.75 7.375 10.03 7.745 ;
  LAYER M4 ;
        RECT 9.725 7.16 10.055 7.96 ;
  LAYER M2 ;
        RECT 1.56 1.12 1.88 1.4 ;
  LAYER M3 ;
        RECT 1.58 1.1 1.86 1.42 ;
  LAYER M2 ;
        RECT 3.28 1.12 3.6 1.4 ;
  LAYER M3 ;
        RECT 3.3 1.1 3.58 1.42 ;
  LAYER M2 ;
        RECT 9.73 7.84 10.05 8.12 ;
  LAYER M3 ;
        RECT 9.75 7.82 10.03 8.14 ;
  LAYER M3 ;
        RECT 3.3 7.375 3.58 7.745 ;
  LAYER M4 ;
        RECT 3.275 7.16 3.605 7.96 ;
  LAYER M3 ;
        RECT 9.75 7.375 10.03 7.745 ;
  LAYER M4 ;
        RECT 9.725 7.16 10.055 7.96 ;
  LAYER M2 ;
        RECT 10.58 7 11.78 7.28 ;
  LAYER M3 ;
        RECT 11.04 8.24 11.32 14.44 ;
  LAYER M2 ;
        RECT 11.02 7 11.34 7.28 ;
  LAYER M3 ;
        RECT 11.04 7.14 11.32 8.4 ;
  LAYER M2 ;
        RECT 11.02 7 11.34 7.28 ;
  LAYER M3 ;
        RECT 11.04 6.98 11.32 7.3 ;
  LAYER M2 ;
        RECT 11.02 7 11.34 7.28 ;
  LAYER M3 ;
        RECT 11.04 6.98 11.32 7.3 ;
  LAYER M2 ;
        RECT 11.44 6.58 12.64 6.86 ;
  LAYER M3 ;
        RECT 12.76 8.24 13.04 14.44 ;
  LAYER M2 ;
        RECT 12.31 6.58 12.63 6.86 ;
  LAYER M3 ;
        RECT 12.33 6.72 12.61 7.56 ;
  LAYER M2 ;
        RECT 12.47 7.42 12.9 7.7 ;
  LAYER M3 ;
        RECT 12.76 7.56 13.04 8.4 ;
  LAYER M2 ;
        RECT 12.31 6.58 12.63 6.86 ;
  LAYER M3 ;
        RECT 12.33 6.56 12.61 6.88 ;
  LAYER M2 ;
        RECT 12.31 7.42 12.63 7.7 ;
  LAYER M3 ;
        RECT 12.33 7.4 12.61 7.72 ;
  LAYER M2 ;
        RECT 12.74 7.42 13.06 7.7 ;
  LAYER M3 ;
        RECT 12.76 7.4 13.04 7.72 ;
  LAYER M2 ;
        RECT 12.31 6.58 12.63 6.86 ;
  LAYER M3 ;
        RECT 12.33 6.56 12.61 6.88 ;
  LAYER M2 ;
        RECT 12.31 7.42 12.63 7.7 ;
  LAYER M3 ;
        RECT 12.33 7.4 12.61 7.72 ;
  LAYER M2 ;
        RECT 12.74 7.42 13.06 7.7 ;
  LAYER M3 ;
        RECT 12.76 7.4 13.04 7.72 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 6.88 ;
  LAYER M3 ;
        RECT 7.6 8.24 7.88 14.44 ;
  LAYER M2 ;
        RECT 14.02 7 15.22 7.28 ;
  LAYER M2 ;
        RECT 14.88 7.84 16.08 8.12 ;
  LAYER M3 ;
        RECT 8.46 6.72 8.74 7.56 ;
  LAYER M2 ;
        RECT 7.74 7.42 8.6 7.7 ;
  LAYER M3 ;
        RECT 7.6 7.56 7.88 8.4 ;
  LAYER M3 ;
        RECT 8.46 6.115 8.74 6.485 ;
  LAYER M4 ;
        RECT 8.6 5.9 13.33 6.7 ;
  LAYER M3 ;
        RECT 13.19 6.3 13.47 7.14 ;
  LAYER M2 ;
        RECT 13.33 7 14.19 7.28 ;
  LAYER M2 ;
        RECT 14.89 7 15.21 7.28 ;
  LAYER M3 ;
        RECT 14.91 7.14 15.19 7.98 ;
  LAYER M2 ;
        RECT 14.89 7.84 15.21 8.12 ;
  LAYER M2 ;
        RECT 7.58 7.42 7.9 7.7 ;
  LAYER M3 ;
        RECT 7.6 7.4 7.88 7.72 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 7.58 7.42 7.9 7.7 ;
  LAYER M3 ;
        RECT 7.6 7.4 7.88 7.72 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 7.58 7.42 7.9 7.7 ;
  LAYER M3 ;
        RECT 7.6 7.4 7.88 7.72 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 13.17 7 13.49 7.28 ;
  LAYER M3 ;
        RECT 13.19 6.98 13.47 7.3 ;
  LAYER M3 ;
        RECT 8.46 6.115 8.74 6.485 ;
  LAYER M4 ;
        RECT 8.435 5.9 8.765 6.7 ;
  LAYER M3 ;
        RECT 13.19 6.115 13.47 6.485 ;
  LAYER M4 ;
        RECT 13.165 5.9 13.495 6.7 ;
  LAYER M2 ;
        RECT 7.58 7.42 7.9 7.7 ;
  LAYER M3 ;
        RECT 7.6 7.4 7.88 7.72 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 13.17 7 13.49 7.28 ;
  LAYER M3 ;
        RECT 13.19 6.98 13.47 7.3 ;
  LAYER M3 ;
        RECT 8.46 6.115 8.74 6.485 ;
  LAYER M4 ;
        RECT 8.435 5.9 8.765 6.7 ;
  LAYER M3 ;
        RECT 13.19 6.115 13.47 6.485 ;
  LAYER M4 ;
        RECT 13.165 5.9 13.495 6.7 ;
  LAYER M2 ;
        RECT 7.58 7.42 7.9 7.7 ;
  LAYER M3 ;
        RECT 7.6 7.4 7.88 7.72 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 13.17 7 13.49 7.28 ;
  LAYER M3 ;
        RECT 13.19 6.98 13.47 7.3 ;
  LAYER M2 ;
        RECT 14.89 7 15.21 7.28 ;
  LAYER M3 ;
        RECT 14.91 6.98 15.19 7.3 ;
  LAYER M2 ;
        RECT 14.89 7.84 15.21 8.12 ;
  LAYER M3 ;
        RECT 14.91 7.82 15.19 8.14 ;
  LAYER M3 ;
        RECT 8.46 6.115 8.74 6.485 ;
  LAYER M4 ;
        RECT 8.435 5.9 8.765 6.7 ;
  LAYER M3 ;
        RECT 13.19 6.115 13.47 6.485 ;
  LAYER M4 ;
        RECT 13.165 5.9 13.495 6.7 ;
  LAYER M2 ;
        RECT 7.58 7.42 7.9 7.7 ;
  LAYER M3 ;
        RECT 7.6 7.4 7.88 7.72 ;
  LAYER M2 ;
        RECT 8.44 7.42 8.76 7.7 ;
  LAYER M3 ;
        RECT 8.46 7.4 8.74 7.72 ;
  LAYER M2 ;
        RECT 13.17 7 13.49 7.28 ;
  LAYER M3 ;
        RECT 13.19 6.98 13.47 7.3 ;
  LAYER M2 ;
        RECT 14.89 7 15.21 7.28 ;
  LAYER M3 ;
        RECT 14.91 6.98 15.19 7.3 ;
  LAYER M2 ;
        RECT 14.89 7.84 15.21 8.12 ;
  LAYER M3 ;
        RECT 14.91 7.82 15.19 8.14 ;
  LAYER M3 ;
        RECT 8.46 6.115 8.74 6.485 ;
  LAYER M4 ;
        RECT 8.435 5.9 8.765 6.7 ;
  LAYER M3 ;
        RECT 13.19 6.115 13.47 6.485 ;
  LAYER M4 ;
        RECT 13.165 5.9 13.495 6.7 ;
  LAYER M1 ;
        RECT 1.165 7.895 1.415 11.425 ;
  LAYER M1 ;
        RECT 1.165 11.675 1.415 12.685 ;
  LAYER M1 ;
        RECT 1.165 13.775 1.415 14.785 ;
  LAYER M1 ;
        RECT 0.735 7.895 0.985 11.425 ;
  LAYER M1 ;
        RECT 1.595 7.895 1.845 11.425 ;
  LAYER M2 ;
        RECT 0.69 8.26 1.89 8.54 ;
  LAYER M2 ;
        RECT 0.69 14.14 1.89 14.42 ;
  LAYER M2 ;
        RECT 0.26 7.84 1.46 8.12 ;
  LAYER M2 ;
        RECT 0.26 12.04 1.46 12.32 ;
  LAYER M3 ;
        RECT 1.58 8.24 1.86 14.44 ;
  LAYER M1 ;
        RECT 1.165 3.695 1.415 7.225 ;
  LAYER M1 ;
        RECT 1.165 2.435 1.415 3.445 ;
  LAYER M1 ;
        RECT 1.165 0.335 1.415 1.345 ;
  LAYER M1 ;
        RECT 0.735 3.695 0.985 7.225 ;
  LAYER M1 ;
        RECT 1.595 3.695 1.845 7.225 ;
  LAYER M2 ;
        RECT 0.69 6.58 1.89 6.86 ;
  LAYER M2 ;
        RECT 0.69 0.7 1.89 0.98 ;
  LAYER M2 ;
        RECT 0.26 7 1.46 7.28 ;
  LAYER M2 ;
        RECT 0.26 2.8 1.46 3.08 ;
  LAYER M3 ;
        RECT 1.58 0.68 1.86 6.88 ;
  LAYER M1 ;
        RECT 11.485 3.695 11.735 7.225 ;
  LAYER M1 ;
        RECT 11.485 2.435 11.735 3.445 ;
  LAYER M1 ;
        RECT 11.485 0.335 11.735 1.345 ;
  LAYER M1 ;
        RECT 11.055 3.695 11.305 7.225 ;
  LAYER M1 ;
        RECT 11.915 3.695 12.165 7.225 ;
  LAYER M1 ;
        RECT 12.345 3.695 12.595 7.225 ;
  LAYER M1 ;
        RECT 12.345 2.435 12.595 3.445 ;
  LAYER M1 ;
        RECT 12.345 0.335 12.595 1.345 ;
  LAYER M1 ;
        RECT 12.775 3.695 13.025 7.225 ;
  LAYER M2 ;
        RECT 11.01 6.16 13.07 6.44 ;
  LAYER M2 ;
        RECT 11.44 0.7 13.07 0.98 ;
  LAYER M2 ;
        RECT 10.58 7 11.78 7.28 ;
  LAYER M2 ;
        RECT 11.44 6.58 12.64 6.86 ;
  LAYER M2 ;
        RECT 10.58 2.8 11.78 3.08 ;
  LAYER M2 ;
        RECT 11.44 2.38 12.64 2.66 ;
  LAYER M3 ;
        RECT 12.76 0.68 13.04 6.46 ;
  LAYER M1 ;
        RECT 14.925 3.695 15.175 7.225 ;
  LAYER M1 ;
        RECT 14.925 2.435 15.175 3.445 ;
  LAYER M1 ;
        RECT 14.925 0.335 15.175 1.345 ;
  LAYER M1 ;
        RECT 14.495 3.695 14.745 7.225 ;
  LAYER M1 ;
        RECT 15.355 3.695 15.605 7.225 ;
  LAYER M2 ;
        RECT 14.45 6.58 15.65 6.86 ;
  LAYER M2 ;
        RECT 14.45 0.7 15.65 0.98 ;
  LAYER M2 ;
        RECT 14.02 7 15.22 7.28 ;
  LAYER M2 ;
        RECT 14.02 2.8 15.22 3.08 ;
  LAYER M3 ;
        RECT 15.34 0.68 15.62 6.88 ;
  LAYER M1 ;
        RECT 15.785 7.895 16.035 11.425 ;
  LAYER M1 ;
        RECT 15.785 11.675 16.035 12.685 ;
  LAYER M1 ;
        RECT 15.785 13.775 16.035 14.785 ;
  LAYER M1 ;
        RECT 15.355 7.895 15.605 11.425 ;
  LAYER M1 ;
        RECT 16.215 7.895 16.465 11.425 ;
  LAYER M2 ;
        RECT 15.31 8.26 16.51 8.54 ;
  LAYER M2 ;
        RECT 15.31 14.14 16.51 14.42 ;
  LAYER M2 ;
        RECT 14.88 7.84 16.08 8.12 ;
  LAYER M2 ;
        RECT 14.88 12.04 16.08 12.32 ;
  LAYER M3 ;
        RECT 16.2 8.24 16.48 14.44 ;
  LAYER M1 ;
        RECT 6.325 3.695 6.575 7.225 ;
  LAYER M1 ;
        RECT 6.325 2.435 6.575 3.445 ;
  LAYER M1 ;
        RECT 6.325 0.335 6.575 1.345 ;
  LAYER M1 ;
        RECT 5.895 3.695 6.145 7.225 ;
  LAYER M1 ;
        RECT 6.755 3.695 7.005 7.225 ;
  LAYER M2 ;
        RECT 5.85 6.58 7.05 6.86 ;
  LAYER M2 ;
        RECT 5.85 0.7 7.05 0.98 ;
  LAYER M2 ;
        RECT 5.42 7 6.62 7.28 ;
  LAYER M2 ;
        RECT 5.42 2.8 6.62 3.08 ;
  LAYER M3 ;
        RECT 6.74 0.68 7.02 6.88 ;
  LAYER M1 ;
        RECT 8.905 3.695 9.155 7.225 ;
  LAYER M1 ;
        RECT 8.905 2.435 9.155 3.445 ;
  LAYER M1 ;
        RECT 8.905 0.335 9.155 1.345 ;
  LAYER M1 ;
        RECT 9.335 3.695 9.585 7.225 ;
  LAYER M1 ;
        RECT 8.475 3.695 8.725 7.225 ;
  LAYER M2 ;
        RECT 8.43 6.58 9.63 6.86 ;
  LAYER M2 ;
        RECT 8.43 0.7 9.63 0.98 ;
  LAYER M2 ;
        RECT 8.86 7 10.06 7.28 ;
  LAYER M2 ;
        RECT 8.86 2.8 10.06 3.08 ;
  LAYER M3 ;
        RECT 8.46 0.68 8.74 6.88 ;
  LAYER M1 ;
        RECT 8.045 7.895 8.295 11.425 ;
  LAYER M1 ;
        RECT 8.045 11.675 8.295 12.685 ;
  LAYER M1 ;
        RECT 8.045 13.775 8.295 14.785 ;
  LAYER M1 ;
        RECT 8.475 7.895 8.725 11.425 ;
  LAYER M1 ;
        RECT 7.615 7.895 7.865 11.425 ;
  LAYER M2 ;
        RECT 7.57 8.26 8.77 8.54 ;
  LAYER M2 ;
        RECT 7.57 14.14 8.77 14.42 ;
  LAYER M2 ;
        RECT 8 7.84 9.2 8.12 ;
  LAYER M2 ;
        RECT 8 12.04 9.2 12.32 ;
  LAYER M3 ;
        RECT 7.6 8.24 7.88 14.44 ;
  LAYER M1 ;
        RECT 3.745 3.695 3.995 7.225 ;
  LAYER M1 ;
        RECT 3.745 2.435 3.995 3.445 ;
  LAYER M1 ;
        RECT 3.745 0.335 3.995 1.345 ;
  LAYER M1 ;
        RECT 4.175 3.695 4.425 7.225 ;
  LAYER M1 ;
        RECT 3.315 3.695 3.565 7.225 ;
  LAYER M2 ;
        RECT 3.27 6.58 4.47 6.86 ;
  LAYER M2 ;
        RECT 3.27 0.7 4.47 0.98 ;
  LAYER M2 ;
        RECT 3.7 7 4.9 7.28 ;
  LAYER M2 ;
        RECT 3.7 2.8 4.9 3.08 ;
  LAYER M3 ;
        RECT 3.3 0.68 3.58 6.88 ;
  LAYER M1 ;
        RECT 10.625 7.895 10.875 11.425 ;
  LAYER M1 ;
        RECT 10.625 11.675 10.875 12.685 ;
  LAYER M1 ;
        RECT 10.625 13.775 10.875 14.785 ;
  LAYER M1 ;
        RECT 10.195 7.895 10.445 11.425 ;
  LAYER M1 ;
        RECT 11.055 7.895 11.305 11.425 ;
  LAYER M2 ;
        RECT 10.15 8.26 11.35 8.54 ;
  LAYER M2 ;
        RECT 10.15 14.14 11.35 14.42 ;
  LAYER M2 ;
        RECT 9.72 7.84 10.92 8.12 ;
  LAYER M2 ;
        RECT 9.72 12.04 10.92 12.32 ;
  LAYER M3 ;
        RECT 11.04 8.24 11.32 14.44 ;
  LAYER M1 ;
        RECT 13.205 7.895 13.455 11.425 ;
  LAYER M1 ;
        RECT 13.205 11.675 13.455 12.685 ;
  LAYER M1 ;
        RECT 13.205 13.775 13.455 14.785 ;
  LAYER M1 ;
        RECT 13.635 7.895 13.885 11.425 ;
  LAYER M1 ;
        RECT 12.775 7.895 13.025 11.425 ;
  LAYER M2 ;
        RECT 12.73 8.26 13.93 8.54 ;
  LAYER M2 ;
        RECT 12.73 14.14 13.93 14.42 ;
  LAYER M2 ;
        RECT 13.16 7.84 14.36 8.12 ;
  LAYER M2 ;
        RECT 13.16 12.04 14.36 12.32 ;
  LAYER M3 ;
        RECT 12.76 8.24 13.04 14.44 ;
  END 
END TEST
