magic
tech sky130A
magscale 1 2
timestamp 1676559991
<< nwell >>
rect 0 0 688 1512
<< pmos >>
rect 200 399 230 735
rect 286 399 316 735
rect 372 399 402 735
rect 458 399 488 735
<< pdiff >>
rect 147 585 200 735
rect 147 551 155 585
rect 189 551 200 585
rect 147 517 200 551
rect 147 483 155 517
rect 189 483 200 517
rect 147 449 200 483
rect 147 415 155 449
rect 189 415 200 449
rect 147 399 200 415
rect 230 585 286 735
rect 230 551 241 585
rect 275 551 286 585
rect 230 517 286 551
rect 230 483 241 517
rect 275 483 286 517
rect 230 449 286 483
rect 230 415 241 449
rect 275 415 286 449
rect 230 399 286 415
rect 316 585 372 735
rect 316 551 327 585
rect 361 551 372 585
rect 316 517 372 551
rect 316 483 327 517
rect 361 483 372 517
rect 316 449 372 483
rect 316 415 327 449
rect 361 415 372 449
rect 316 399 372 415
rect 402 585 458 735
rect 402 551 413 585
rect 447 551 458 585
rect 402 517 458 551
rect 402 483 413 517
rect 447 483 458 517
rect 402 449 458 483
rect 402 415 413 449
rect 447 415 458 449
rect 402 399 458 415
rect 488 585 541 735
rect 488 551 499 585
rect 533 551 541 585
rect 488 517 541 551
rect 488 483 499 517
rect 533 483 541 517
rect 488 449 541 483
rect 488 415 499 449
rect 533 415 541 449
rect 488 399 541 415
<< pdiffc >>
rect 155 551 189 585
rect 155 483 189 517
rect 155 415 189 449
rect 241 551 275 585
rect 241 483 275 517
rect 241 415 275 449
rect 327 551 361 585
rect 327 483 361 517
rect 327 415 361 449
rect 413 551 447 585
rect 413 483 447 517
rect 413 415 447 449
rect 499 551 533 585
rect 499 483 533 517
rect 499 415 533 449
<< nsubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
rect 413 1361 447 1456
rect 413 1232 447 1327
<< nsubdiffcont >>
rect 241 1327 275 1361
rect 413 1327 447 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 735 230 897
rect 286 735 316 897
rect 372 941 488 951
rect 372 907 413 941
rect 447 907 488 941
rect 372 897 488 907
rect 372 735 402 897
rect 458 735 488 897
rect 200 252 230 399
rect 286 252 316 399
rect 372 252 402 399
rect 458 252 488 399
<< polycont >>
rect 241 907 275 941
rect 413 907 447 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 405 1361 455 1445
rect 405 1327 413 1361
rect 447 1327 455 1361
rect 405 1243 455 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 405 991 413 1025
rect 447 991 455 1025
rect 405 941 455 991
rect 405 907 413 941
rect 447 907 455 941
rect 405 823 455 907
rect 147 585 197 773
rect 147 551 155 585
rect 189 551 197 585
rect 147 517 197 551
rect 147 483 155 517
rect 189 483 197 517
rect 147 449 197 483
rect 147 415 155 449
rect 189 415 197 449
rect 147 269 197 415
rect 147 235 155 269
rect 189 235 197 269
rect 147 67 197 235
rect 233 585 283 773
rect 233 551 241 585
rect 275 551 283 585
rect 233 517 283 551
rect 233 483 241 517
rect 275 483 283 517
rect 233 449 283 483
rect 233 415 241 449
rect 275 415 283 449
rect 233 101 283 415
rect 233 67 241 101
rect 275 67 283 101
rect 319 585 369 773
rect 319 551 327 585
rect 361 551 369 585
rect 319 517 369 551
rect 319 483 327 517
rect 361 483 369 517
rect 319 449 369 483
rect 319 415 327 449
rect 361 415 369 449
rect 319 269 369 415
rect 319 235 327 269
rect 361 235 369 269
rect 319 67 369 235
rect 405 585 455 773
rect 405 551 413 585
rect 447 551 455 585
rect 405 517 455 551
rect 405 483 413 517
rect 447 483 455 517
rect 405 449 455 483
rect 405 415 413 449
rect 447 415 455 449
rect 405 185 455 415
rect 405 151 413 185
rect 447 151 455 185
rect 405 67 455 151
rect 491 585 541 773
rect 491 551 499 585
rect 533 551 541 585
rect 491 517 541 551
rect 491 483 499 517
rect 533 483 541 517
rect 491 449 541 483
rect 491 415 499 449
rect 533 415 541 449
rect 491 269 541 415
rect 491 235 499 269
rect 533 235 541 269
rect 491 67 541 235
<< viali >>
rect 241 1327 275 1361
rect 413 1327 447 1361
rect 241 907 275 941
rect 413 991 447 1025
rect 155 235 189 269
rect 241 67 275 101
rect 327 235 361 269
rect 413 151 447 185
rect 499 235 533 269
<< metal1 >>
rect 224 1370 550 1372
rect 224 1361 490 1370
rect 224 1327 241 1361
rect 275 1327 413 1361
rect 447 1327 490 1361
rect 224 1318 490 1327
rect 542 1318 550 1370
rect 224 1316 550 1318
rect 224 1025 464 1036
rect 224 991 413 1025
rect 447 991 464 1025
rect 224 980 464 991
rect 52 941 292 952
rect 52 907 241 941
rect 275 907 292 941
rect 52 896 292 907
rect 138 278 550 280
rect 138 269 490 278
rect 138 235 155 269
rect 189 235 327 269
rect 361 235 490 269
rect 138 226 490 235
rect 542 226 550 278
rect 138 224 550 226
rect 224 185 464 196
rect 224 151 413 185
rect 447 151 464 185
rect 224 140 464 151
rect 52 101 292 112
rect 52 67 241 101
rect 275 67 292 101
rect 52 56 292 67
<< via1 >>
rect 490 1318 542 1370
rect 490 269 542 278
rect 490 235 499 269
rect 499 235 533 269
rect 533 235 542 269
rect 490 226 542 235
<< metal2 >>
rect 488 1370 544 1376
rect 488 1318 490 1370
rect 542 1318 544 1370
rect 488 278 544 1318
rect 488 226 490 278
rect 542 226 544 278
rect 488 220 544 226
<< end >>
