magic
tech sky130A
magscale 1 2
timestamp 1677523798
<< error_s >>
rect -2546 3750 -2488 3756
rect -2546 3716 -2534 3750
rect -2546 3710 -2488 3716
rect -2642 3454 -2584 3460
rect -2642 3420 -2630 3454
rect -2642 3414 -2584 3420
rect -2100 3282 -2048 3888
rect -1644 3872 -1574 3888
rect -1818 3750 -1760 3756
rect -1818 3716 -1806 3750
rect -1818 3710 -1760 3716
rect -1914 3454 -1856 3460
rect -1914 3420 -1902 3454
rect -1914 3414 -1856 3420
rect -1390 3282 -1320 3872
rect -1108 3734 -1050 3740
rect -1108 3700 -1096 3734
rect -1108 3694 -1050 3700
rect -1204 3438 -1146 3444
rect -1204 3404 -1192 3438
rect -1204 3398 -1146 3404
rect -1786 3116 -1728 3122
rect -1786 3082 -1774 3116
rect -1786 3076 -1728 3082
rect -1026 3066 -968 3072
rect -2530 3050 -2472 3056
rect -2530 3016 -2518 3050
rect -1026 3032 -1014 3066
rect -1026 3026 -968 3032
rect -2530 3010 -2472 3016
rect -1882 2922 -1824 2928
rect -1882 2888 -1870 2922
rect -1882 2882 -1824 2888
rect -1122 2872 -1064 2878
rect -2626 2856 -2568 2862
rect -2626 2822 -2614 2856
rect -1122 2838 -1110 2872
rect -1122 2832 -1064 2838
rect -2626 2816 -2568 2822
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC1
timestamp 1677523798
transform 1 0 6024 0 1 3322
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC2
timestamp 1677523798
transform 1 0 6080 0 1 -3052
box -3186 -3040 3186 3040
use sky130_fd_pr__cap_mim_m3_1_3HBNLG  XC3
timestamp 1677523798
transform 1 0 -548 0 1 -3084
box -3186 -3040 3186 3040
use sky130_fd_pr__pfet_01v8_MQKFPY  XM1
timestamp 1677523798
transform 1 0 -1837 0 1 3585
box -263 -303 263 303
use sky130_fd_pr__pfet_01v8_MQKFPY  XM2
timestamp 1677523798
transform 1 0 -2565 0 1 3585
box -263 -303 263 303
use sky130_fd_pr__pfet_01v8_MQKFPY  XM3
timestamp 1677523798
transform 1 0 -1127 0 1 3569
box -263 -303 263 303
use sky130_fd_pr__nfet_01v8_MVW3GX  XM4
timestamp 1677523798
transform 1 0 -2549 0 1 2936
box -263 -252 263 252
use sky130_fd_pr__nfet_01v8_MVW3GX  XM5
timestamp 1677523798
transform 1 0 -1805 0 1 3002
box -263 -252 263 252
use sky130_fd_pr__nfet_01v8_MVW3GX  XM6
timestamp 1677523798
transform 1 0 -1045 0 1 2952
box -263 -252 263 252
<< end >>
