magic
tech sky130A
magscale 1 2
timestamp 1676559991
<< pwell >>
rect 215 1206 301 1482
rect 121 457 395 677
<< nmos >>
rect 200 483 230 651
rect 286 483 316 651
<< ndiff >>
rect 147 601 200 651
rect 147 567 155 601
rect 189 567 200 601
rect 147 533 200 567
rect 147 499 155 533
rect 189 499 200 533
rect 147 483 200 499
rect 230 601 286 651
rect 230 567 241 601
rect 275 567 286 601
rect 230 533 286 567
rect 230 499 241 533
rect 275 499 286 533
rect 230 483 286 499
rect 316 601 369 651
rect 316 567 327 601
rect 361 567 369 601
rect 316 533 369 567
rect 316 499 327 533
rect 361 499 369 533
rect 316 483 369 499
<< ndiffc >>
rect 155 567 189 601
rect 155 499 189 533
rect 241 567 275 601
rect 241 499 275 533
rect 327 567 361 601
rect 327 499 361 533
<< psubdiff >>
rect 241 1361 275 1456
rect 241 1232 275 1327
<< psubdiffcont >>
rect 241 1327 275 1361
<< poly >>
rect 200 941 316 951
rect 200 907 241 941
rect 275 907 316 941
rect 200 897 316 907
rect 200 651 230 897
rect 286 651 316 897
rect 200 252 230 483
rect 286 252 316 483
<< polycont >>
rect 241 907 275 941
<< locali >>
rect 233 1361 283 1445
rect 233 1327 241 1361
rect 275 1327 283 1361
rect 233 1243 283 1327
rect 233 941 283 1025
rect 233 907 241 941
rect 275 907 283 941
rect 233 823 283 907
rect 147 601 197 773
rect 147 567 155 601
rect 189 567 197 601
rect 147 533 197 567
rect 147 499 155 533
rect 189 499 197 533
rect 147 185 197 499
rect 147 151 155 185
rect 189 151 197 185
rect 147 67 197 151
rect 233 601 283 773
rect 233 567 241 601
rect 275 567 283 601
rect 233 533 283 567
rect 233 499 241 533
rect 275 499 283 533
rect 233 101 283 499
rect 233 67 241 101
rect 275 67 283 101
rect 319 601 369 773
rect 319 567 327 601
rect 361 567 369 601
rect 319 533 369 567
rect 319 499 327 533
rect 361 499 369 533
rect 319 185 369 499
rect 319 151 327 185
rect 361 151 369 185
rect 319 67 369 151
<< viali >>
rect 241 1327 275 1361
rect 241 907 275 941
rect 155 151 189 185
rect 241 67 275 101
rect 327 151 361 185
<< metal1 >>
rect 138 1370 378 1372
rect 138 1361 318 1370
rect 138 1327 241 1361
rect 275 1327 318 1361
rect 138 1318 318 1327
rect 370 1318 378 1370
rect 138 1316 378 1318
rect 52 941 292 952
rect 52 907 241 941
rect 275 907 292 941
rect 52 896 292 907
rect 138 194 378 196
rect 138 185 318 194
rect 138 151 155 185
rect 189 151 318 185
rect 138 142 318 151
rect 370 142 378 194
rect 138 140 378 142
rect 52 101 292 112
rect 52 67 241 101
rect 275 67 292 101
rect 52 56 292 67
<< via1 >>
rect 318 1318 370 1370
rect 318 185 370 194
rect 318 151 327 185
rect 327 151 361 185
rect 361 151 370 185
rect 318 142 370 151
<< metal2 >>
rect 316 1370 372 1376
rect 316 1318 318 1370
rect 370 1318 372 1370
rect 316 194 372 1318
rect 316 142 318 194
rect 370 142 372 194
rect 316 136 372 142
<< end >>
